`timescale 1ns / 1ps

module tb_motion_estimation;

    // ==========================================
    // 1. 訊號宣告
    // ==========================================
    reg clk;
    reg rst_n;
    reg start;
    wire done;
    wire [15:0] min_sad;
    wire signed [5:0] mv_x; // 假設 Range +/- 31 以內
    wire signed [5:0] mv_y;

    // 定義記憶體來存放 Python 產生的資料
    reg [7:0] cur_mem [0:255];          // 16x16 = 256 pixels
    reg [7:0] ref_window_mem [0:1023];  // Search Window (假設夠大)

    // ==========================================
    // 2. 讀取 Python 檔案 ($readmemh)
    // ==========================================
    initial begin
        $display("Loading Hex files generated by Python...");
        // 讀取 cur_block.hex 到 cur_mem
        $readmemh("cur_block.hex", cur_mem);
        // 讀取 search_window.hex 到 ref_window_mem
        $readmemh("search_window.hex", ref_window_mem);
        $display("Data loaded successfully.");
    end

    // ==========================================
    // 3. 實例化你的設計 (DUT - Device Under Test)
    // ==========================================
    // 注意：這裡假設你有一個叫做 hexagon_me_top 的模組
    // 你需要根據論文去實作這個模組
    /*
    hexagon_me_top u_dut (
        .clk(clk),
        .rst_n(rst_n),
        .start(start),
        // 這裡需要透過記憶體介面把資料傳進去，或者直接在內部讀取 mem
        .current_pixel_in(...), 
        .done(done),
        .final_mv_x(mv_x),
        .final_mv_y(mv_y),
        .final_sad(min_sad)
    );
    */

    // ==========================================
    // 4. 時脈產生 (Clock Generation)
    // ==========================================
    initial clk = 0;
    always #5 clk = ~clk; // 100MHz (10ns period)

    // ==========================================
    // 5. 測試流程控制
    // ==========================================
    initial begin
        // 初始化訊號
        rst_n = 0;
        start = 0;
        
        // Reset 釋放
        #100;
        rst_n = 1;
        
        // 啟動運算
        #20;
        start = 1;
        #10;
        start = 0;

        // 等待完成 (模擬等待)
        // 實際情況要偵測 done 訊號
        wait(done == 1); 
        
        // 顯示結果
        $display("----------------------------------");
        $display("Simulation Done!");
        $display("HW Output MV: (%d, %d)", mv_x, mv_y);
        $display("HW Output SAD: %d", min_sad);
        $display("----------------------------------");
        
        // 也可以把結果寫回文字檔讓 Python 讀
        // $fdisplay(...);

        $finish;
    end

    // 安全機制：跑太久就強制停止
    initial begin
        #100000; 
        $display("Timeout! Simulation took too long.");
        $finish;
    end

endmodule