magic
tech sky130A
magscale 1 2
timestamp 1766521404
<< obsli1 >>
rect 1104 2159 156400 157233
<< obsm1 >>
rect 14 1708 157214 157264
<< metal2 >>
rect 18 158919 74 159719
rect 2594 158919 2650 159719
rect 5814 158919 5870 159719
rect 9034 158919 9090 159719
rect 12254 158919 12310 159719
rect 15474 158919 15530 159719
rect 18050 158919 18106 159719
rect 21270 158919 21326 159719
rect 24490 158919 24546 159719
rect 27710 158919 27766 159719
rect 30930 158919 30986 159719
rect 33506 158919 33562 159719
rect 36726 158919 36782 159719
rect 39946 158919 40002 159719
rect 43166 158919 43222 159719
rect 46386 158919 46442 159719
rect 48962 158919 49018 159719
rect 52182 158919 52238 159719
rect 55402 158919 55458 159719
rect 58622 158919 58678 159719
rect 61842 158919 61898 159719
rect 64418 158919 64474 159719
rect 67638 158919 67694 159719
rect 70858 158919 70914 159719
rect 74078 158919 74134 159719
rect 77298 158919 77354 159719
rect 79874 158919 79930 159719
rect 83094 158919 83150 159719
rect 86314 158919 86370 159719
rect 89534 158919 89590 159719
rect 92754 158919 92810 159719
rect 95330 158919 95386 159719
rect 98550 158919 98606 159719
rect 101770 158919 101826 159719
rect 104990 158919 105046 159719
rect 108210 158919 108266 159719
rect 110786 158919 110842 159719
rect 114006 158919 114062 159719
rect 117226 158919 117282 159719
rect 120446 158919 120502 159719
rect 123666 158919 123722 159719
rect 126242 158919 126298 159719
rect 129462 158919 129518 159719
rect 132682 158919 132738 159719
rect 135902 158919 135958 159719
rect 139122 158919 139178 159719
rect 141698 158919 141754 159719
rect 144918 158919 144974 159719
rect 148138 158919 148194 159719
rect 151358 158919 151414 159719
rect 154578 158919 154634 159719
rect 157154 158919 157210 159719
rect 18 0 74 800
rect 2594 0 2650 800
rect 5814 0 5870 800
rect 9034 0 9090 800
rect 12254 0 12310 800
rect 15474 0 15530 800
rect 18050 0 18106 800
rect 21270 0 21326 800
rect 24490 0 24546 800
rect 27710 0 27766 800
rect 30930 0 30986 800
rect 33506 0 33562 800
rect 36726 0 36782 800
rect 39946 0 40002 800
rect 43166 0 43222 800
rect 46386 0 46442 800
rect 48962 0 49018 800
rect 52182 0 52238 800
rect 55402 0 55458 800
rect 58622 0 58678 800
rect 61842 0 61898 800
rect 64418 0 64474 800
rect 67638 0 67694 800
rect 70858 0 70914 800
rect 74078 0 74134 800
rect 77298 0 77354 800
rect 79874 0 79930 800
rect 83094 0 83150 800
rect 86314 0 86370 800
rect 89534 0 89590 800
rect 92754 0 92810 800
rect 95330 0 95386 800
rect 98550 0 98606 800
rect 101770 0 101826 800
rect 104990 0 105046 800
rect 108210 0 108266 800
rect 110786 0 110842 800
rect 114006 0 114062 800
rect 117226 0 117282 800
rect 120446 0 120502 800
rect 123666 0 123722 800
rect 126242 0 126298 800
rect 129462 0 129518 800
rect 132682 0 132738 800
rect 135902 0 135958 800
rect 139122 0 139178 800
rect 141698 0 141754 800
rect 144918 0 144974 800
rect 148138 0 148194 800
rect 151358 0 151414 800
rect 154578 0 154634 800
rect 157154 0 157210 800
<< obsm2 >>
rect 130 158863 2538 159066
rect 2706 158863 5758 159066
rect 5926 158863 8978 159066
rect 9146 158863 12198 159066
rect 12366 158863 15418 159066
rect 15586 158863 17994 159066
rect 18162 158863 21214 159066
rect 21382 158863 24434 159066
rect 24602 158863 27654 159066
rect 27822 158863 30874 159066
rect 31042 158863 33450 159066
rect 33618 158863 36670 159066
rect 36838 158863 39890 159066
rect 40058 158863 43110 159066
rect 43278 158863 46330 159066
rect 46498 158863 48906 159066
rect 49074 158863 52126 159066
rect 52294 158863 55346 159066
rect 55514 158863 58566 159066
rect 58734 158863 61786 159066
rect 61954 158863 64362 159066
rect 64530 158863 67582 159066
rect 67750 158863 70802 159066
rect 70970 158863 74022 159066
rect 74190 158863 77242 159066
rect 77410 158863 79818 159066
rect 79986 158863 83038 159066
rect 83206 158863 86258 159066
rect 86426 158863 89478 159066
rect 89646 158863 92698 159066
rect 92866 158863 95274 159066
rect 95442 158863 98494 159066
rect 98662 158863 101714 159066
rect 101882 158863 104934 159066
rect 105102 158863 108154 159066
rect 108322 158863 110730 159066
rect 110898 158863 113950 159066
rect 114118 158863 117170 159066
rect 117338 158863 120390 159066
rect 120558 158863 123610 159066
rect 123778 158863 126186 159066
rect 126354 158863 129406 159066
rect 129574 158863 132626 159066
rect 132794 158863 135846 159066
rect 136014 158863 139066 159066
rect 139234 158863 141642 159066
rect 141810 158863 144862 159066
rect 145030 158863 148082 159066
rect 148250 158863 151302 159066
rect 151470 158863 154522 159066
rect 154690 158863 157098 159066
rect 20 856 157208 158863
rect 130 734 2538 856
rect 2706 734 5758 856
rect 5926 734 8978 856
rect 9146 734 12198 856
rect 12366 734 15418 856
rect 15586 734 17994 856
rect 18162 734 21214 856
rect 21382 734 24434 856
rect 24602 734 27654 856
rect 27822 734 30874 856
rect 31042 734 33450 856
rect 33618 734 36670 856
rect 36838 734 39890 856
rect 40058 734 43110 856
rect 43278 734 46330 856
rect 46498 734 48906 856
rect 49074 734 52126 856
rect 52294 734 55346 856
rect 55514 734 58566 856
rect 58734 734 61786 856
rect 61954 734 64362 856
rect 64530 734 67582 856
rect 67750 734 70802 856
rect 70970 734 74022 856
rect 74190 734 77242 856
rect 77410 734 79818 856
rect 79986 734 83038 856
rect 83206 734 86258 856
rect 86426 734 89478 856
rect 89646 734 92698 856
rect 92866 734 95274 856
rect 95442 734 98494 856
rect 98662 734 101714 856
rect 101882 734 104934 856
rect 105102 734 108154 856
rect 108322 734 110730 856
rect 110898 734 113950 856
rect 114118 734 117170 856
rect 117338 734 120390 856
rect 120558 734 123610 856
rect 123778 734 126186 856
rect 126354 734 129406 856
rect 129574 734 132626 856
rect 132794 734 135846 856
rect 136014 734 139066 856
rect 139234 734 141642 856
rect 141810 734 144862 856
rect 145030 734 148082 856
rect 148250 734 151302 856
rect 151470 734 154522 856
rect 154690 734 157098 856
<< metal3 >>
rect 0 156408 800 156528
rect 156775 156408 157575 156528
rect 0 153008 800 153128
rect 156775 153008 157575 153128
rect 0 149608 800 149728
rect 156775 149608 157575 149728
rect 0 146208 800 146328
rect 156775 146208 157575 146328
rect 0 143488 800 143608
rect 156775 143488 157575 143608
rect 0 140088 800 140208
rect 156775 140088 157575 140208
rect 0 136688 800 136808
rect 156775 136688 157575 136808
rect 0 133288 800 133408
rect 156775 133288 157575 133408
rect 0 129888 800 130008
rect 156775 129888 157575 130008
rect 0 127168 800 127288
rect 156775 127168 157575 127288
rect 0 123768 800 123888
rect 156775 123768 157575 123888
rect 0 120368 800 120488
rect 156775 120368 157575 120488
rect 0 116968 800 117088
rect 156775 116968 157575 117088
rect 0 113568 800 113688
rect 156775 113568 157575 113688
rect 0 110848 800 110968
rect 156775 110848 157575 110968
rect 0 107448 800 107568
rect 156775 107448 157575 107568
rect 0 104048 800 104168
rect 156775 104048 157575 104168
rect 0 100648 800 100768
rect 156775 100648 157575 100768
rect 0 97248 800 97368
rect 156775 97248 157575 97368
rect 0 94528 800 94648
rect 156775 94528 157575 94648
rect 0 91128 800 91248
rect 156775 91128 157575 91248
rect 0 87728 800 87848
rect 156775 87728 157575 87848
rect 0 84328 800 84448
rect 156775 84328 157575 84448
rect 0 80928 800 81048
rect 156775 80928 157575 81048
rect 0 78208 800 78328
rect 156775 78208 157575 78328
rect 0 74808 800 74928
rect 156775 74808 157575 74928
rect 0 71408 800 71528
rect 156775 71408 157575 71528
rect 0 68008 800 68128
rect 156775 68008 157575 68128
rect 0 64608 800 64728
rect 156775 64608 157575 64728
rect 0 61888 800 62008
rect 156775 61888 157575 62008
rect 0 58488 800 58608
rect 156775 58488 157575 58608
rect 0 55088 800 55208
rect 156775 55088 157575 55208
rect 0 51688 800 51808
rect 156775 51688 157575 51808
rect 0 48288 800 48408
rect 156775 48288 157575 48408
rect 0 45568 800 45688
rect 156775 45568 157575 45688
rect 0 42168 800 42288
rect 156775 42168 157575 42288
rect 0 38768 800 38888
rect 156775 38768 157575 38888
rect 0 35368 800 35488
rect 156775 35368 157575 35488
rect 0 31968 800 32088
rect 156775 31968 157575 32088
rect 0 29248 800 29368
rect 156775 29248 157575 29368
rect 0 25848 800 25968
rect 156775 25848 157575 25968
rect 0 22448 800 22568
rect 156775 22448 157575 22568
rect 0 19048 800 19168
rect 156775 19048 157575 19168
rect 0 15648 800 15768
rect 156775 15648 157575 15768
rect 0 12928 800 13048
rect 156775 12928 157575 13048
rect 0 9528 800 9648
rect 156775 9528 157575 9648
rect 0 6128 800 6248
rect 156775 6128 157575 6248
rect 0 2728 800 2848
rect 156775 2728 157575 2848
<< obsm3 >>
rect 798 156608 156775 157249
rect 880 156328 156695 156608
rect 798 153208 156775 156328
rect 880 152928 156695 153208
rect 798 149808 156775 152928
rect 880 149528 156695 149808
rect 798 146408 156775 149528
rect 880 146128 156695 146408
rect 798 143688 156775 146128
rect 880 143408 156695 143688
rect 798 140288 156775 143408
rect 880 140008 156695 140288
rect 798 136888 156775 140008
rect 880 136608 156695 136888
rect 798 133488 156775 136608
rect 880 133208 156695 133488
rect 798 130088 156775 133208
rect 880 129808 156695 130088
rect 798 127368 156775 129808
rect 880 127088 156695 127368
rect 798 123968 156775 127088
rect 880 123688 156695 123968
rect 798 120568 156775 123688
rect 880 120288 156695 120568
rect 798 117168 156775 120288
rect 880 116888 156695 117168
rect 798 113768 156775 116888
rect 880 113488 156695 113768
rect 798 111048 156775 113488
rect 880 110768 156695 111048
rect 798 107648 156775 110768
rect 880 107368 156695 107648
rect 798 104248 156775 107368
rect 880 103968 156695 104248
rect 798 100848 156775 103968
rect 880 100568 156695 100848
rect 798 97448 156775 100568
rect 880 97168 156695 97448
rect 798 94728 156775 97168
rect 880 94448 156695 94728
rect 798 91328 156775 94448
rect 880 91048 156695 91328
rect 798 87928 156775 91048
rect 880 87648 156695 87928
rect 798 84528 156775 87648
rect 880 84248 156695 84528
rect 798 81128 156775 84248
rect 880 80848 156695 81128
rect 798 78408 156775 80848
rect 880 78128 156695 78408
rect 798 75008 156775 78128
rect 880 74728 156695 75008
rect 798 71608 156775 74728
rect 880 71328 156695 71608
rect 798 68208 156775 71328
rect 880 67928 156695 68208
rect 798 64808 156775 67928
rect 880 64528 156695 64808
rect 798 62088 156775 64528
rect 880 61808 156695 62088
rect 798 58688 156775 61808
rect 880 58408 156695 58688
rect 798 55288 156775 58408
rect 880 55008 156695 55288
rect 798 51888 156775 55008
rect 880 51608 156695 51888
rect 798 48488 156775 51608
rect 880 48208 156695 48488
rect 798 45768 156775 48208
rect 880 45488 156695 45768
rect 798 42368 156775 45488
rect 880 42088 156695 42368
rect 798 38968 156775 42088
rect 880 38688 156695 38968
rect 798 35568 156775 38688
rect 880 35288 156695 35568
rect 798 32168 156775 35288
rect 880 31888 156695 32168
rect 798 29448 156775 31888
rect 880 29168 156695 29448
rect 798 26048 156775 29168
rect 880 25768 156695 26048
rect 798 22648 156775 25768
rect 880 22368 156695 22648
rect 798 19248 156775 22368
rect 880 18968 156695 19248
rect 798 15848 156775 18968
rect 880 15568 156695 15848
rect 798 13128 156775 15568
rect 880 12848 156695 13128
rect 798 9728 156775 12848
rect 880 9448 156695 9728
rect 798 6328 156775 9448
rect 880 6048 156695 6328
rect 798 2928 156775 6048
rect 880 2648 156695 2928
rect 798 2143 156775 2648
<< metal4 >>
rect 4208 2128 4528 157264
rect 4868 2128 5188 157264
rect 34928 2128 35248 157264
rect 35588 2128 35908 157264
rect 65648 2128 65968 157264
rect 66308 2128 66628 157264
rect 96368 2128 96688 157264
rect 97028 2128 97348 157264
rect 127088 2128 127408 157264
rect 127748 2128 128068 157264
<< obsm4 >>
rect 5395 2619 34848 153237
rect 35328 2619 35508 153237
rect 35988 2619 65568 153237
rect 66048 2619 66228 153237
rect 66708 2619 96288 153237
rect 96768 2619 96948 153237
rect 97428 2619 127008 153237
rect 127488 2619 127668 153237
rect 128148 2619 153581 153237
<< metal5 >>
rect 1056 128550 156448 128870
rect 1056 127890 156448 128210
rect 1056 97914 156448 98234
rect 1056 97254 156448 97574
rect 1056 67278 156448 67598
rect 1056 66618 156448 66938
rect 1056 36642 156448 36962
rect 1056 35982 156448 36302
rect 1056 6006 156448 6326
rect 1056 5346 156448 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 157264 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 157264 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 157264 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 97028 2128 97348 157264 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127748 2128 128068 157264 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 156448 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 156448 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 67278 156448 67598 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 97914 156448 98234 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 128550 156448 128870 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 157264 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157264 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157264 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157264 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 157264 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 156448 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 156448 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66618 156448 66938 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 97254 156448 97574 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 127890 156448 128210 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 15474 0 15530 800 6 clk
port 3 nsew signal input
rlabel metal2 s 64418 158919 64474 159719 6 done
port 4 nsew signal output
rlabel metal2 s 52182 158919 52238 159719 6 frame_start_addr[0]
port 5 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 frame_start_addr[10]
port 6 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 frame_start_addr[11]
port 7 nsew signal input
rlabel metal3 s 156775 29248 157575 29368 6 frame_start_addr[12]
port 8 nsew signal input
rlabel metal3 s 0 149608 800 149728 6 frame_start_addr[13]
port 9 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 frame_start_addr[14]
port 10 nsew signal input
rlabel metal3 s 156775 9528 157575 9648 6 frame_start_addr[15]
port 11 nsew signal input
rlabel metal2 s 33506 158919 33562 159719 6 frame_start_addr[16]
port 12 nsew signal input
rlabel metal3 s 156775 87728 157575 87848 6 frame_start_addr[17]
port 13 nsew signal input
rlabel metal3 s 156775 120368 157575 120488 6 frame_start_addr[18]
port 14 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 frame_start_addr[19]
port 15 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 frame_start_addr[1]
port 16 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 frame_start_addr[20]
port 17 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 frame_start_addr[21]
port 18 nsew signal input
rlabel metal2 s 98550 158919 98606 159719 6 frame_start_addr[22]
port 19 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 frame_start_addr[23]
port 20 nsew signal input
rlabel metal2 s 154578 158919 154634 159719 6 frame_start_addr[24]
port 21 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 frame_start_addr[25]
port 22 nsew signal input
rlabel metal2 s 48962 158919 49018 159719 6 frame_start_addr[26]
port 23 nsew signal input
rlabel metal3 s 156775 45568 157575 45688 6 frame_start_addr[27]
port 24 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 frame_start_addr[28]
port 25 nsew signal input
rlabel metal3 s 156775 84328 157575 84448 6 frame_start_addr[29]
port 26 nsew signal input
rlabel metal2 s 30930 158919 30986 159719 6 frame_start_addr[2]
port 27 nsew signal input
rlabel metal2 s 9034 158919 9090 159719 6 frame_start_addr[30]
port 28 nsew signal input
rlabel metal2 s 129462 158919 129518 159719 6 frame_start_addr[31]
port 29 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 frame_start_addr[3]
port 30 nsew signal input
rlabel metal3 s 156775 143488 157575 143608 6 frame_start_addr[4]
port 31 nsew signal input
rlabel metal3 s 156775 123768 157575 123888 6 frame_start_addr[5]
port 32 nsew signal input
rlabel metal3 s 156775 64608 157575 64728 6 frame_start_addr[6]
port 33 nsew signal input
rlabel metal3 s 156775 51688 157575 51808 6 frame_start_addr[7]
port 34 nsew signal input
rlabel metal2 s 58622 158919 58678 159719 6 frame_start_addr[8]
port 35 nsew signal input
rlabel metal2 s 77298 158919 77354 159719 6 frame_start_addr[9]
port 36 nsew signal input
rlabel metal2 s 139122 158919 139178 159719 6 mb_x_pos[0]
port 37 nsew signal input
rlabel metal3 s 156775 19048 157575 19168 6 mb_x_pos[10]
port 38 nsew signal input
rlabel metal2 s 117226 158919 117282 159719 6 mb_x_pos[11]
port 39 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 mb_x_pos[12]
port 40 nsew signal input
rlabel metal2 s 135902 158919 135958 159719 6 mb_x_pos[13]
port 41 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 mb_x_pos[14]
port 42 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 mb_x_pos[15]
port 43 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 mb_x_pos[16]
port 44 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 mb_x_pos[17]
port 45 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 mb_x_pos[18]
port 46 nsew signal input
rlabel metal3 s 156775 80928 157575 81048 6 mb_x_pos[19]
port 47 nsew signal input
rlabel metal3 s 156775 153008 157575 153128 6 mb_x_pos[1]
port 48 nsew signal input
rlabel metal2 s 123666 158919 123722 159719 6 mb_x_pos[20]
port 49 nsew signal input
rlabel metal2 s 18 158919 74 159719 6 mb_x_pos[21]
port 50 nsew signal input
rlabel metal2 s 61842 158919 61898 159719 6 mb_x_pos[22]
port 51 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 mb_x_pos[23]
port 52 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 mb_x_pos[24]
port 53 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 mb_x_pos[25]
port 54 nsew signal input
rlabel metal3 s 156775 42168 157575 42288 6 mb_x_pos[26]
port 55 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 mb_x_pos[27]
port 56 nsew signal input
rlabel metal3 s 156775 129888 157575 130008 6 mb_x_pos[28]
port 57 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 mb_x_pos[29]
port 58 nsew signal input
rlabel metal2 s 36726 158919 36782 159719 6 mb_x_pos[2]
port 59 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 mb_x_pos[30]
port 60 nsew signal input
rlabel metal2 s 43166 158919 43222 159719 6 mb_x_pos[31]
port 61 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 mb_x_pos[3]
port 62 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 mb_x_pos[4]
port 63 nsew signal input
rlabel metal2 s 46386 158919 46442 159719 6 mb_x_pos[5]
port 64 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 mb_x_pos[6]
port 65 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 mb_x_pos[7]
port 66 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 mb_x_pos[8]
port 67 nsew signal input
rlabel metal3 s 156775 2728 157575 2848 6 mb_x_pos[9]
port 68 nsew signal input
rlabel metal3 s 156775 94528 157575 94648 6 mb_y_pos[0]
port 69 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 mb_y_pos[10]
port 70 nsew signal input
rlabel metal2 s 114006 158919 114062 159719 6 mb_y_pos[11]
port 71 nsew signal input
rlabel metal2 s 39946 158919 40002 159719 6 mb_y_pos[12]
port 72 nsew signal input
rlabel metal3 s 156775 156408 157575 156528 6 mb_y_pos[13]
port 73 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 mb_y_pos[14]
port 74 nsew signal input
rlabel metal3 s 0 120368 800 120488 6 mb_y_pos[15]
port 75 nsew signal input
rlabel metal3 s 156775 97248 157575 97368 6 mb_y_pos[16]
port 76 nsew signal input
rlabel metal3 s 156775 136688 157575 136808 6 mb_y_pos[17]
port 77 nsew signal input
rlabel metal3 s 156775 35368 157575 35488 6 mb_y_pos[18]
port 78 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 mb_y_pos[19]
port 79 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 mb_y_pos[1]
port 80 nsew signal input
rlabel metal3 s 156775 25848 157575 25968 6 mb_y_pos[20]
port 81 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 mb_y_pos[21]
port 82 nsew signal input
rlabel metal3 s 156775 55088 157575 55208 6 mb_y_pos[22]
port 83 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 mb_y_pos[23]
port 84 nsew signal input
rlabel metal3 s 156775 91128 157575 91248 6 mb_y_pos[24]
port 85 nsew signal input
rlabel metal2 s 157154 158919 157210 159719 6 mb_y_pos[25]
port 86 nsew signal input
rlabel metal2 s 120446 158919 120502 159719 6 mb_y_pos[26]
port 87 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 mb_y_pos[27]
port 88 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 mb_y_pos[28]
port 89 nsew signal input
rlabel metal3 s 0 143488 800 143608 6 mb_y_pos[29]
port 90 nsew signal input
rlabel metal2 s 89534 158919 89590 159719 6 mb_y_pos[2]
port 91 nsew signal input
rlabel metal2 s 132682 158919 132738 159719 6 mb_y_pos[30]
port 92 nsew signal input
rlabel metal2 s 21270 158919 21326 159719 6 mb_y_pos[31]
port 93 nsew signal input
rlabel metal2 s 67638 158919 67694 159719 6 mb_y_pos[3]
port 94 nsew signal input
rlabel metal3 s 156775 113568 157575 113688 6 mb_y_pos[4]
port 95 nsew signal input
rlabel metal2 s 86314 158919 86370 159719 6 mb_y_pos[5]
port 96 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 mb_y_pos[6]
port 97 nsew signal input
rlabel metal3 s 156775 127168 157575 127288 6 mb_y_pos[7]
port 98 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 mb_y_pos[8]
port 99 nsew signal input
rlabel metal2 s 18050 158919 18106 159719 6 mb_y_pos[9]
port 100 nsew signal input
rlabel metal3 s 156775 104048 157575 104168 6 mem_addr[0]
port 101 nsew signal output
rlabel metal3 s 156775 146208 157575 146328 6 mem_addr[10]
port 102 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 mem_addr[11]
port 103 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 mem_addr[12]
port 104 nsew signal output
rlabel metal2 s 5814 158919 5870 159719 6 mem_addr[13]
port 105 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 mem_addr[14]
port 106 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 mem_addr[15]
port 107 nsew signal output
rlabel metal3 s 156775 12928 157575 13048 6 mem_addr[16]
port 108 nsew signal output
rlabel metal3 s 0 146208 800 146328 6 mem_addr[17]
port 109 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 mem_addr[18]
port 110 nsew signal output
rlabel metal2 s 95330 158919 95386 159719 6 mem_addr[19]
port 111 nsew signal output
rlabel metal2 s 101770 158919 101826 159719 6 mem_addr[1]
port 112 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 mem_addr[20]
port 113 nsew signal output
rlabel metal2 s 83094 158919 83150 159719 6 mem_addr[21]
port 114 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 mem_addr[22]
port 115 nsew signal output
rlabel metal2 s 148138 158919 148194 159719 6 mem_addr[23]
port 116 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 mem_addr[24]
port 117 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 mem_addr[25]
port 118 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 mem_addr[26]
port 119 nsew signal output
rlabel metal3 s 156775 22448 157575 22568 6 mem_addr[27]
port 120 nsew signal output
rlabel metal3 s 156775 68008 157575 68128 6 mem_addr[28]
port 121 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 mem_addr[29]
port 122 nsew signal output
rlabel metal3 s 156775 100648 157575 100768 6 mem_addr[2]
port 123 nsew signal output
rlabel metal3 s 156775 6128 157575 6248 6 mem_addr[30]
port 124 nsew signal output
rlabel metal2 s 12254 158919 12310 159719 6 mem_addr[31]
port 125 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 mem_addr[3]
port 126 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 mem_addr[4]
port 127 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 mem_addr[5]
port 128 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 mem_addr[6]
port 129 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 mem_addr[7]
port 130 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 mem_addr[8]
port 131 nsew signal output
rlabel metal2 s 141698 158919 141754 159719 6 mem_addr[9]
port 132 nsew signal output
rlabel metal3 s 156775 71408 157575 71528 6 mem_rdata[0]
port 133 nsew signal input
rlabel metal2 s 55402 158919 55458 159719 6 mem_rdata[1]
port 134 nsew signal input
rlabel metal2 s 79874 158919 79930 159719 6 mem_rdata[2]
port 135 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 mem_rdata[3]
port 136 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 mem_rdata[4]
port 137 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 mem_rdata[5]
port 138 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 mem_rdata[6]
port 139 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 mem_rdata[7]
port 140 nsew signal input
rlabel metal3 s 156775 140088 157575 140208 6 mv_x[0]
port 141 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 mv_x[1]
port 142 nsew signal output
rlabel metal2 s 92754 158919 92810 159719 6 mv_x[2]
port 143 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 mv_x[3]
port 144 nsew signal output
rlabel metal3 s 156775 48288 157575 48408 6 mv_x[4]
port 145 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 mv_x[5]
port 146 nsew signal output
rlabel metal2 s 27710 158919 27766 159719 6 mv_y[0]
port 147 nsew signal output
rlabel metal3 s 156775 78208 157575 78328 6 mv_y[1]
port 148 nsew signal output
rlabel metal3 s 0 153008 800 153128 6 mv_y[2]
port 149 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 mv_y[3]
port 150 nsew signal output
rlabel metal3 s 156775 133288 157575 133408 6 mv_y[4]
port 151 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 mv_y[5]
port 152 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 ref_start_addr[0]
port 153 nsew signal input
rlabel metal3 s 156775 58488 157575 58608 6 ref_start_addr[10]
port 154 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 ref_start_addr[11]
port 155 nsew signal input
rlabel metal3 s 156775 15648 157575 15768 6 ref_start_addr[12]
port 156 nsew signal input
rlabel metal2 s 2594 158919 2650 159719 6 ref_start_addr[13]
port 157 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 ref_start_addr[14]
port 158 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 ref_start_addr[15]
port 159 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 ref_start_addr[16]
port 160 nsew signal input
rlabel metal3 s 156775 38768 157575 38888 6 ref_start_addr[17]
port 161 nsew signal input
rlabel metal3 s 156775 149608 157575 149728 6 ref_start_addr[18]
port 162 nsew signal input
rlabel metal3 s 156775 107448 157575 107568 6 ref_start_addr[19]
port 163 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 ref_start_addr[1]
port 164 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 ref_start_addr[20]
port 165 nsew signal input
rlabel metal3 s 156775 61888 157575 62008 6 ref_start_addr[21]
port 166 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 ref_start_addr[22]
port 167 nsew signal input
rlabel metal3 s 156775 116968 157575 117088 6 ref_start_addr[23]
port 168 nsew signal input
rlabel metal2 s 151358 158919 151414 159719 6 ref_start_addr[24]
port 169 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 ref_start_addr[25]
port 170 nsew signal input
rlabel metal2 s 144918 158919 144974 159719 6 ref_start_addr[26]
port 171 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 ref_start_addr[27]
port 172 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 ref_start_addr[28]
port 173 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 ref_start_addr[29]
port 174 nsew signal input
rlabel metal2 s 18 0 74 800 6 ref_start_addr[2]
port 175 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 ref_start_addr[30]
port 176 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 ref_start_addr[31]
port 177 nsew signal input
rlabel metal2 s 15474 158919 15530 159719 6 ref_start_addr[3]
port 178 nsew signal input
rlabel metal2 s 74078 158919 74134 159719 6 ref_start_addr[4]
port 179 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 ref_start_addr[5]
port 180 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 ref_start_addr[6]
port 181 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 ref_start_addr[7]
port 182 nsew signal input
rlabel metal2 s 104990 158919 105046 159719 6 ref_start_addr[8]
port 183 nsew signal input
rlabel metal2 s 70858 158919 70914 159719 6 ref_start_addr[9]
port 184 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 rst_n
port 185 nsew signal input
rlabel metal2 s 126242 158919 126298 159719 6 sad[0]
port 186 nsew signal output
rlabel metal3 s 156775 31968 157575 32088 6 sad[10]
port 187 nsew signal output
rlabel metal3 s 0 127168 800 127288 6 sad[11]
port 188 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 sad[12]
port 189 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 sad[13]
port 190 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 sad[14]
port 191 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 sad[15]
port 192 nsew signal output
rlabel metal3 s 156775 110848 157575 110968 6 sad[1]
port 193 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 sad[2]
port 194 nsew signal output
rlabel metal2 s 110786 158919 110842 159719 6 sad[3]
port 195 nsew signal output
rlabel metal2 s 108210 158919 108266 159719 6 sad[4]
port 196 nsew signal output
rlabel metal3 s 0 156408 800 156528 6 sad[5]
port 197 nsew signal output
rlabel metal2 s 24490 158919 24546 159719 6 sad[6]
port 198 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 sad[7]
port 199 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 sad[8]
port 200 nsew signal output
rlabel metal3 s 0 136688 800 136808 6 sad[9]
port 201 nsew signal output
rlabel metal3 s 156775 74808 157575 74928 6 start
port 202 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 157575 159719
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 41648364
string GDS_FILE /openlane/designs/hexbs/runs/RUN_2025.12.23_20.06.50/results/signoff/hexbs_top.magic.gds
string GDS_START 1263198
<< end >>

