module hexbs_top (clk,
    done,
    rst_n,
    start,
    frame_start_addr,
    mb_x_pos,
    mb_y_pos,
    mem_addr,
    mem_rdata,
    mv_x,
    mv_y,
    ref_start_addr,
    sad);
 input clk;
 output done;
 input rst_n;
 input start;
 input [31:0] frame_start_addr;
 input [31:0] mb_x_pos;
 input [31:0] mb_y_pos;
 output [31:0] mem_addr;
 input [7:0] mem_rdata;
 output [5:0] mv_x;
 output [5:0] mv_y;
 input [31:0] ref_start_addr;
 output [15:0] sad;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire \best_cand_x[0] ;
 wire \best_cand_x[1] ;
 wire \best_cand_x[2] ;
 wire \best_cand_x[3] ;
 wire \best_cand_x[4] ;
 wire \best_cand_x[5] ;
 wire \best_cand_x[6] ;
 wire \best_cand_y[0] ;
 wire \best_cand_y[1] ;
 wire \best_cand_y[2] ;
 wire \best_cand_y[3] ;
 wire \best_cand_y[4] ;
 wire \best_cand_y[5] ;
 wire \best_cand_y[6] ;
 wire \best_point_idx[0] ;
 wire \best_point_idx[1] ;
 wire \best_point_idx[2] ;
 wire \best_point_idx[3] ;
 wire \cand_x[0] ;
 wire \cand_x[1] ;
 wire \cand_x[2] ;
 wire \cand_x[3] ;
 wire \cand_x[4] ;
 wire \cand_x[5] ;
 wire \cand_x[6] ;
 wire \cand_y[0] ;
 wire \cand_y[1] ;
 wire \cand_y[2] ;
 wire \cand_y[3] ;
 wire \cand_y[4] ;
 wire \cand_y[5] ;
 wire \cand_y[6] ;
 wire \center_x[0] ;
 wire \center_x[1] ;
 wire \center_x[2] ;
 wire \center_x[3] ;
 wire \center_x[4] ;
 wire \center_x[5] ;
 wire \center_x[6] ;
 wire \center_y[0] ;
 wire \center_y[1] ;
 wire \center_y[2] ;
 wire \center_y[3] ;
 wire \center_y[4] ;
 wire \center_y[5] ;
 wire \center_y[6] ;
 wire \cur_mb_mem[0][0] ;
 wire \cur_mb_mem[0][1] ;
 wire \cur_mb_mem[0][2] ;
 wire \cur_mb_mem[0][3] ;
 wire \cur_mb_mem[0][4] ;
 wire \cur_mb_mem[0][5] ;
 wire \cur_mb_mem[0][6] ;
 wire \cur_mb_mem[0][7] ;
 wire \cur_mb_mem[100][0] ;
 wire \cur_mb_mem[100][1] ;
 wire \cur_mb_mem[100][2] ;
 wire \cur_mb_mem[100][3] ;
 wire \cur_mb_mem[100][4] ;
 wire \cur_mb_mem[100][5] ;
 wire \cur_mb_mem[100][6] ;
 wire \cur_mb_mem[100][7] ;
 wire \cur_mb_mem[101][0] ;
 wire \cur_mb_mem[101][1] ;
 wire \cur_mb_mem[101][2] ;
 wire \cur_mb_mem[101][3] ;
 wire \cur_mb_mem[101][4] ;
 wire \cur_mb_mem[101][5] ;
 wire \cur_mb_mem[101][6] ;
 wire \cur_mb_mem[101][7] ;
 wire \cur_mb_mem[102][0] ;
 wire \cur_mb_mem[102][1] ;
 wire \cur_mb_mem[102][2] ;
 wire \cur_mb_mem[102][3] ;
 wire \cur_mb_mem[102][4] ;
 wire \cur_mb_mem[102][5] ;
 wire \cur_mb_mem[102][6] ;
 wire \cur_mb_mem[102][7] ;
 wire \cur_mb_mem[103][0] ;
 wire \cur_mb_mem[103][1] ;
 wire \cur_mb_mem[103][2] ;
 wire \cur_mb_mem[103][3] ;
 wire \cur_mb_mem[103][4] ;
 wire \cur_mb_mem[103][5] ;
 wire \cur_mb_mem[103][6] ;
 wire \cur_mb_mem[103][7] ;
 wire \cur_mb_mem[104][0] ;
 wire \cur_mb_mem[104][1] ;
 wire \cur_mb_mem[104][2] ;
 wire \cur_mb_mem[104][3] ;
 wire \cur_mb_mem[104][4] ;
 wire \cur_mb_mem[104][5] ;
 wire \cur_mb_mem[104][6] ;
 wire \cur_mb_mem[104][7] ;
 wire \cur_mb_mem[105][0] ;
 wire \cur_mb_mem[105][1] ;
 wire \cur_mb_mem[105][2] ;
 wire \cur_mb_mem[105][3] ;
 wire \cur_mb_mem[105][4] ;
 wire \cur_mb_mem[105][5] ;
 wire \cur_mb_mem[105][6] ;
 wire \cur_mb_mem[105][7] ;
 wire \cur_mb_mem[106][0] ;
 wire \cur_mb_mem[106][1] ;
 wire \cur_mb_mem[106][2] ;
 wire \cur_mb_mem[106][3] ;
 wire \cur_mb_mem[106][4] ;
 wire \cur_mb_mem[106][5] ;
 wire \cur_mb_mem[106][6] ;
 wire \cur_mb_mem[106][7] ;
 wire \cur_mb_mem[107][0] ;
 wire \cur_mb_mem[107][1] ;
 wire \cur_mb_mem[107][2] ;
 wire \cur_mb_mem[107][3] ;
 wire \cur_mb_mem[107][4] ;
 wire \cur_mb_mem[107][5] ;
 wire \cur_mb_mem[107][6] ;
 wire \cur_mb_mem[107][7] ;
 wire \cur_mb_mem[108][0] ;
 wire \cur_mb_mem[108][1] ;
 wire \cur_mb_mem[108][2] ;
 wire \cur_mb_mem[108][3] ;
 wire \cur_mb_mem[108][4] ;
 wire \cur_mb_mem[108][5] ;
 wire \cur_mb_mem[108][6] ;
 wire \cur_mb_mem[108][7] ;
 wire \cur_mb_mem[109][0] ;
 wire \cur_mb_mem[109][1] ;
 wire \cur_mb_mem[109][2] ;
 wire \cur_mb_mem[109][3] ;
 wire \cur_mb_mem[109][4] ;
 wire \cur_mb_mem[109][5] ;
 wire \cur_mb_mem[109][6] ;
 wire \cur_mb_mem[109][7] ;
 wire \cur_mb_mem[10][0] ;
 wire \cur_mb_mem[10][1] ;
 wire \cur_mb_mem[10][2] ;
 wire \cur_mb_mem[10][3] ;
 wire \cur_mb_mem[10][4] ;
 wire \cur_mb_mem[10][5] ;
 wire \cur_mb_mem[10][6] ;
 wire \cur_mb_mem[10][7] ;
 wire \cur_mb_mem[110][0] ;
 wire \cur_mb_mem[110][1] ;
 wire \cur_mb_mem[110][2] ;
 wire \cur_mb_mem[110][3] ;
 wire \cur_mb_mem[110][4] ;
 wire \cur_mb_mem[110][5] ;
 wire \cur_mb_mem[110][6] ;
 wire \cur_mb_mem[110][7] ;
 wire \cur_mb_mem[111][0] ;
 wire \cur_mb_mem[111][1] ;
 wire \cur_mb_mem[111][2] ;
 wire \cur_mb_mem[111][3] ;
 wire \cur_mb_mem[111][4] ;
 wire \cur_mb_mem[111][5] ;
 wire \cur_mb_mem[111][6] ;
 wire \cur_mb_mem[111][7] ;
 wire \cur_mb_mem[112][0] ;
 wire \cur_mb_mem[112][1] ;
 wire \cur_mb_mem[112][2] ;
 wire \cur_mb_mem[112][3] ;
 wire \cur_mb_mem[112][4] ;
 wire \cur_mb_mem[112][5] ;
 wire \cur_mb_mem[112][6] ;
 wire \cur_mb_mem[112][7] ;
 wire \cur_mb_mem[113][0] ;
 wire \cur_mb_mem[113][1] ;
 wire \cur_mb_mem[113][2] ;
 wire \cur_mb_mem[113][3] ;
 wire \cur_mb_mem[113][4] ;
 wire \cur_mb_mem[113][5] ;
 wire \cur_mb_mem[113][6] ;
 wire \cur_mb_mem[113][7] ;
 wire \cur_mb_mem[114][0] ;
 wire \cur_mb_mem[114][1] ;
 wire \cur_mb_mem[114][2] ;
 wire \cur_mb_mem[114][3] ;
 wire \cur_mb_mem[114][4] ;
 wire \cur_mb_mem[114][5] ;
 wire \cur_mb_mem[114][6] ;
 wire \cur_mb_mem[114][7] ;
 wire \cur_mb_mem[115][0] ;
 wire \cur_mb_mem[115][1] ;
 wire \cur_mb_mem[115][2] ;
 wire \cur_mb_mem[115][3] ;
 wire \cur_mb_mem[115][4] ;
 wire \cur_mb_mem[115][5] ;
 wire \cur_mb_mem[115][6] ;
 wire \cur_mb_mem[115][7] ;
 wire \cur_mb_mem[116][0] ;
 wire \cur_mb_mem[116][1] ;
 wire \cur_mb_mem[116][2] ;
 wire \cur_mb_mem[116][3] ;
 wire \cur_mb_mem[116][4] ;
 wire \cur_mb_mem[116][5] ;
 wire \cur_mb_mem[116][6] ;
 wire \cur_mb_mem[116][7] ;
 wire \cur_mb_mem[117][0] ;
 wire \cur_mb_mem[117][1] ;
 wire \cur_mb_mem[117][2] ;
 wire \cur_mb_mem[117][3] ;
 wire \cur_mb_mem[117][4] ;
 wire \cur_mb_mem[117][5] ;
 wire \cur_mb_mem[117][6] ;
 wire \cur_mb_mem[117][7] ;
 wire \cur_mb_mem[118][0] ;
 wire \cur_mb_mem[118][1] ;
 wire \cur_mb_mem[118][2] ;
 wire \cur_mb_mem[118][3] ;
 wire \cur_mb_mem[118][4] ;
 wire \cur_mb_mem[118][5] ;
 wire \cur_mb_mem[118][6] ;
 wire \cur_mb_mem[118][7] ;
 wire \cur_mb_mem[119][0] ;
 wire \cur_mb_mem[119][1] ;
 wire \cur_mb_mem[119][2] ;
 wire \cur_mb_mem[119][3] ;
 wire \cur_mb_mem[119][4] ;
 wire \cur_mb_mem[119][5] ;
 wire \cur_mb_mem[119][6] ;
 wire \cur_mb_mem[119][7] ;
 wire \cur_mb_mem[11][0] ;
 wire \cur_mb_mem[11][1] ;
 wire \cur_mb_mem[11][2] ;
 wire \cur_mb_mem[11][3] ;
 wire \cur_mb_mem[11][4] ;
 wire \cur_mb_mem[11][5] ;
 wire \cur_mb_mem[11][6] ;
 wire \cur_mb_mem[11][7] ;
 wire \cur_mb_mem[120][0] ;
 wire \cur_mb_mem[120][1] ;
 wire \cur_mb_mem[120][2] ;
 wire \cur_mb_mem[120][3] ;
 wire \cur_mb_mem[120][4] ;
 wire \cur_mb_mem[120][5] ;
 wire \cur_mb_mem[120][6] ;
 wire \cur_mb_mem[120][7] ;
 wire \cur_mb_mem[121][0] ;
 wire \cur_mb_mem[121][1] ;
 wire \cur_mb_mem[121][2] ;
 wire \cur_mb_mem[121][3] ;
 wire \cur_mb_mem[121][4] ;
 wire \cur_mb_mem[121][5] ;
 wire \cur_mb_mem[121][6] ;
 wire \cur_mb_mem[121][7] ;
 wire \cur_mb_mem[122][0] ;
 wire \cur_mb_mem[122][1] ;
 wire \cur_mb_mem[122][2] ;
 wire \cur_mb_mem[122][3] ;
 wire \cur_mb_mem[122][4] ;
 wire \cur_mb_mem[122][5] ;
 wire \cur_mb_mem[122][6] ;
 wire \cur_mb_mem[122][7] ;
 wire \cur_mb_mem[123][0] ;
 wire \cur_mb_mem[123][1] ;
 wire \cur_mb_mem[123][2] ;
 wire \cur_mb_mem[123][3] ;
 wire \cur_mb_mem[123][4] ;
 wire \cur_mb_mem[123][5] ;
 wire \cur_mb_mem[123][6] ;
 wire \cur_mb_mem[123][7] ;
 wire \cur_mb_mem[124][0] ;
 wire \cur_mb_mem[124][1] ;
 wire \cur_mb_mem[124][2] ;
 wire \cur_mb_mem[124][3] ;
 wire \cur_mb_mem[124][4] ;
 wire \cur_mb_mem[124][5] ;
 wire \cur_mb_mem[124][6] ;
 wire \cur_mb_mem[124][7] ;
 wire \cur_mb_mem[125][0] ;
 wire \cur_mb_mem[125][1] ;
 wire \cur_mb_mem[125][2] ;
 wire \cur_mb_mem[125][3] ;
 wire \cur_mb_mem[125][4] ;
 wire \cur_mb_mem[125][5] ;
 wire \cur_mb_mem[125][6] ;
 wire \cur_mb_mem[125][7] ;
 wire \cur_mb_mem[126][0] ;
 wire \cur_mb_mem[126][1] ;
 wire \cur_mb_mem[126][2] ;
 wire \cur_mb_mem[126][3] ;
 wire \cur_mb_mem[126][4] ;
 wire \cur_mb_mem[126][5] ;
 wire \cur_mb_mem[126][6] ;
 wire \cur_mb_mem[126][7] ;
 wire \cur_mb_mem[127][0] ;
 wire \cur_mb_mem[127][1] ;
 wire \cur_mb_mem[127][2] ;
 wire \cur_mb_mem[127][3] ;
 wire \cur_mb_mem[127][4] ;
 wire \cur_mb_mem[127][5] ;
 wire \cur_mb_mem[127][6] ;
 wire \cur_mb_mem[127][7] ;
 wire \cur_mb_mem[128][0] ;
 wire \cur_mb_mem[128][1] ;
 wire \cur_mb_mem[128][2] ;
 wire \cur_mb_mem[128][3] ;
 wire \cur_mb_mem[128][4] ;
 wire \cur_mb_mem[128][5] ;
 wire \cur_mb_mem[128][6] ;
 wire \cur_mb_mem[128][7] ;
 wire \cur_mb_mem[129][0] ;
 wire \cur_mb_mem[129][1] ;
 wire \cur_mb_mem[129][2] ;
 wire \cur_mb_mem[129][3] ;
 wire \cur_mb_mem[129][4] ;
 wire \cur_mb_mem[129][5] ;
 wire \cur_mb_mem[129][6] ;
 wire \cur_mb_mem[129][7] ;
 wire \cur_mb_mem[12][0] ;
 wire \cur_mb_mem[12][1] ;
 wire \cur_mb_mem[12][2] ;
 wire \cur_mb_mem[12][3] ;
 wire \cur_mb_mem[12][4] ;
 wire \cur_mb_mem[12][5] ;
 wire \cur_mb_mem[12][6] ;
 wire \cur_mb_mem[12][7] ;
 wire \cur_mb_mem[130][0] ;
 wire \cur_mb_mem[130][1] ;
 wire \cur_mb_mem[130][2] ;
 wire \cur_mb_mem[130][3] ;
 wire \cur_mb_mem[130][4] ;
 wire \cur_mb_mem[130][5] ;
 wire \cur_mb_mem[130][6] ;
 wire \cur_mb_mem[130][7] ;
 wire \cur_mb_mem[131][0] ;
 wire \cur_mb_mem[131][1] ;
 wire \cur_mb_mem[131][2] ;
 wire \cur_mb_mem[131][3] ;
 wire \cur_mb_mem[131][4] ;
 wire \cur_mb_mem[131][5] ;
 wire \cur_mb_mem[131][6] ;
 wire \cur_mb_mem[131][7] ;
 wire \cur_mb_mem[132][0] ;
 wire \cur_mb_mem[132][1] ;
 wire \cur_mb_mem[132][2] ;
 wire \cur_mb_mem[132][3] ;
 wire \cur_mb_mem[132][4] ;
 wire \cur_mb_mem[132][5] ;
 wire \cur_mb_mem[132][6] ;
 wire \cur_mb_mem[132][7] ;
 wire \cur_mb_mem[133][0] ;
 wire \cur_mb_mem[133][1] ;
 wire \cur_mb_mem[133][2] ;
 wire \cur_mb_mem[133][3] ;
 wire \cur_mb_mem[133][4] ;
 wire \cur_mb_mem[133][5] ;
 wire \cur_mb_mem[133][6] ;
 wire \cur_mb_mem[133][7] ;
 wire \cur_mb_mem[134][0] ;
 wire \cur_mb_mem[134][1] ;
 wire \cur_mb_mem[134][2] ;
 wire \cur_mb_mem[134][3] ;
 wire \cur_mb_mem[134][4] ;
 wire \cur_mb_mem[134][5] ;
 wire \cur_mb_mem[134][6] ;
 wire \cur_mb_mem[134][7] ;
 wire \cur_mb_mem[135][0] ;
 wire \cur_mb_mem[135][1] ;
 wire \cur_mb_mem[135][2] ;
 wire \cur_mb_mem[135][3] ;
 wire \cur_mb_mem[135][4] ;
 wire \cur_mb_mem[135][5] ;
 wire \cur_mb_mem[135][6] ;
 wire \cur_mb_mem[135][7] ;
 wire \cur_mb_mem[136][0] ;
 wire \cur_mb_mem[136][1] ;
 wire \cur_mb_mem[136][2] ;
 wire \cur_mb_mem[136][3] ;
 wire \cur_mb_mem[136][4] ;
 wire \cur_mb_mem[136][5] ;
 wire \cur_mb_mem[136][6] ;
 wire \cur_mb_mem[136][7] ;
 wire \cur_mb_mem[137][0] ;
 wire \cur_mb_mem[137][1] ;
 wire \cur_mb_mem[137][2] ;
 wire \cur_mb_mem[137][3] ;
 wire \cur_mb_mem[137][4] ;
 wire \cur_mb_mem[137][5] ;
 wire \cur_mb_mem[137][6] ;
 wire \cur_mb_mem[137][7] ;
 wire \cur_mb_mem[138][0] ;
 wire \cur_mb_mem[138][1] ;
 wire \cur_mb_mem[138][2] ;
 wire \cur_mb_mem[138][3] ;
 wire \cur_mb_mem[138][4] ;
 wire \cur_mb_mem[138][5] ;
 wire \cur_mb_mem[138][6] ;
 wire \cur_mb_mem[138][7] ;
 wire \cur_mb_mem[139][0] ;
 wire \cur_mb_mem[139][1] ;
 wire \cur_mb_mem[139][2] ;
 wire \cur_mb_mem[139][3] ;
 wire \cur_mb_mem[139][4] ;
 wire \cur_mb_mem[139][5] ;
 wire \cur_mb_mem[139][6] ;
 wire \cur_mb_mem[139][7] ;
 wire \cur_mb_mem[13][0] ;
 wire \cur_mb_mem[13][1] ;
 wire \cur_mb_mem[13][2] ;
 wire \cur_mb_mem[13][3] ;
 wire \cur_mb_mem[13][4] ;
 wire \cur_mb_mem[13][5] ;
 wire \cur_mb_mem[13][6] ;
 wire \cur_mb_mem[13][7] ;
 wire \cur_mb_mem[140][0] ;
 wire \cur_mb_mem[140][1] ;
 wire \cur_mb_mem[140][2] ;
 wire \cur_mb_mem[140][3] ;
 wire \cur_mb_mem[140][4] ;
 wire \cur_mb_mem[140][5] ;
 wire \cur_mb_mem[140][6] ;
 wire \cur_mb_mem[140][7] ;
 wire \cur_mb_mem[141][0] ;
 wire \cur_mb_mem[141][1] ;
 wire \cur_mb_mem[141][2] ;
 wire \cur_mb_mem[141][3] ;
 wire \cur_mb_mem[141][4] ;
 wire \cur_mb_mem[141][5] ;
 wire \cur_mb_mem[141][6] ;
 wire \cur_mb_mem[141][7] ;
 wire \cur_mb_mem[142][0] ;
 wire \cur_mb_mem[142][1] ;
 wire \cur_mb_mem[142][2] ;
 wire \cur_mb_mem[142][3] ;
 wire \cur_mb_mem[142][4] ;
 wire \cur_mb_mem[142][5] ;
 wire \cur_mb_mem[142][6] ;
 wire \cur_mb_mem[142][7] ;
 wire \cur_mb_mem[143][0] ;
 wire \cur_mb_mem[143][1] ;
 wire \cur_mb_mem[143][2] ;
 wire \cur_mb_mem[143][3] ;
 wire \cur_mb_mem[143][4] ;
 wire \cur_mb_mem[143][5] ;
 wire \cur_mb_mem[143][6] ;
 wire \cur_mb_mem[143][7] ;
 wire \cur_mb_mem[144][0] ;
 wire \cur_mb_mem[144][1] ;
 wire \cur_mb_mem[144][2] ;
 wire \cur_mb_mem[144][3] ;
 wire \cur_mb_mem[144][4] ;
 wire \cur_mb_mem[144][5] ;
 wire \cur_mb_mem[144][6] ;
 wire \cur_mb_mem[144][7] ;
 wire \cur_mb_mem[145][0] ;
 wire \cur_mb_mem[145][1] ;
 wire \cur_mb_mem[145][2] ;
 wire \cur_mb_mem[145][3] ;
 wire \cur_mb_mem[145][4] ;
 wire \cur_mb_mem[145][5] ;
 wire \cur_mb_mem[145][6] ;
 wire \cur_mb_mem[145][7] ;
 wire \cur_mb_mem[146][0] ;
 wire \cur_mb_mem[146][1] ;
 wire \cur_mb_mem[146][2] ;
 wire \cur_mb_mem[146][3] ;
 wire \cur_mb_mem[146][4] ;
 wire \cur_mb_mem[146][5] ;
 wire \cur_mb_mem[146][6] ;
 wire \cur_mb_mem[146][7] ;
 wire \cur_mb_mem[147][0] ;
 wire \cur_mb_mem[147][1] ;
 wire \cur_mb_mem[147][2] ;
 wire \cur_mb_mem[147][3] ;
 wire \cur_mb_mem[147][4] ;
 wire \cur_mb_mem[147][5] ;
 wire \cur_mb_mem[147][6] ;
 wire \cur_mb_mem[147][7] ;
 wire \cur_mb_mem[148][0] ;
 wire \cur_mb_mem[148][1] ;
 wire \cur_mb_mem[148][2] ;
 wire \cur_mb_mem[148][3] ;
 wire \cur_mb_mem[148][4] ;
 wire \cur_mb_mem[148][5] ;
 wire \cur_mb_mem[148][6] ;
 wire \cur_mb_mem[148][7] ;
 wire \cur_mb_mem[149][0] ;
 wire \cur_mb_mem[149][1] ;
 wire \cur_mb_mem[149][2] ;
 wire \cur_mb_mem[149][3] ;
 wire \cur_mb_mem[149][4] ;
 wire \cur_mb_mem[149][5] ;
 wire \cur_mb_mem[149][6] ;
 wire \cur_mb_mem[149][7] ;
 wire \cur_mb_mem[14][0] ;
 wire \cur_mb_mem[14][1] ;
 wire \cur_mb_mem[14][2] ;
 wire \cur_mb_mem[14][3] ;
 wire \cur_mb_mem[14][4] ;
 wire \cur_mb_mem[14][5] ;
 wire \cur_mb_mem[14][6] ;
 wire \cur_mb_mem[14][7] ;
 wire \cur_mb_mem[150][0] ;
 wire \cur_mb_mem[150][1] ;
 wire \cur_mb_mem[150][2] ;
 wire \cur_mb_mem[150][3] ;
 wire \cur_mb_mem[150][4] ;
 wire \cur_mb_mem[150][5] ;
 wire \cur_mb_mem[150][6] ;
 wire \cur_mb_mem[150][7] ;
 wire \cur_mb_mem[151][0] ;
 wire \cur_mb_mem[151][1] ;
 wire \cur_mb_mem[151][2] ;
 wire \cur_mb_mem[151][3] ;
 wire \cur_mb_mem[151][4] ;
 wire \cur_mb_mem[151][5] ;
 wire \cur_mb_mem[151][6] ;
 wire \cur_mb_mem[151][7] ;
 wire \cur_mb_mem[152][0] ;
 wire \cur_mb_mem[152][1] ;
 wire \cur_mb_mem[152][2] ;
 wire \cur_mb_mem[152][3] ;
 wire \cur_mb_mem[152][4] ;
 wire \cur_mb_mem[152][5] ;
 wire \cur_mb_mem[152][6] ;
 wire \cur_mb_mem[152][7] ;
 wire \cur_mb_mem[153][0] ;
 wire \cur_mb_mem[153][1] ;
 wire \cur_mb_mem[153][2] ;
 wire \cur_mb_mem[153][3] ;
 wire \cur_mb_mem[153][4] ;
 wire \cur_mb_mem[153][5] ;
 wire \cur_mb_mem[153][6] ;
 wire \cur_mb_mem[153][7] ;
 wire \cur_mb_mem[154][0] ;
 wire \cur_mb_mem[154][1] ;
 wire \cur_mb_mem[154][2] ;
 wire \cur_mb_mem[154][3] ;
 wire \cur_mb_mem[154][4] ;
 wire \cur_mb_mem[154][5] ;
 wire \cur_mb_mem[154][6] ;
 wire \cur_mb_mem[154][7] ;
 wire \cur_mb_mem[155][0] ;
 wire \cur_mb_mem[155][1] ;
 wire \cur_mb_mem[155][2] ;
 wire \cur_mb_mem[155][3] ;
 wire \cur_mb_mem[155][4] ;
 wire \cur_mb_mem[155][5] ;
 wire \cur_mb_mem[155][6] ;
 wire \cur_mb_mem[155][7] ;
 wire \cur_mb_mem[156][0] ;
 wire \cur_mb_mem[156][1] ;
 wire \cur_mb_mem[156][2] ;
 wire \cur_mb_mem[156][3] ;
 wire \cur_mb_mem[156][4] ;
 wire \cur_mb_mem[156][5] ;
 wire \cur_mb_mem[156][6] ;
 wire \cur_mb_mem[156][7] ;
 wire \cur_mb_mem[157][0] ;
 wire \cur_mb_mem[157][1] ;
 wire \cur_mb_mem[157][2] ;
 wire \cur_mb_mem[157][3] ;
 wire \cur_mb_mem[157][4] ;
 wire \cur_mb_mem[157][5] ;
 wire \cur_mb_mem[157][6] ;
 wire \cur_mb_mem[157][7] ;
 wire \cur_mb_mem[158][0] ;
 wire \cur_mb_mem[158][1] ;
 wire \cur_mb_mem[158][2] ;
 wire \cur_mb_mem[158][3] ;
 wire \cur_mb_mem[158][4] ;
 wire \cur_mb_mem[158][5] ;
 wire \cur_mb_mem[158][6] ;
 wire \cur_mb_mem[158][7] ;
 wire \cur_mb_mem[159][0] ;
 wire \cur_mb_mem[159][1] ;
 wire \cur_mb_mem[159][2] ;
 wire \cur_mb_mem[159][3] ;
 wire \cur_mb_mem[159][4] ;
 wire \cur_mb_mem[159][5] ;
 wire \cur_mb_mem[159][6] ;
 wire \cur_mb_mem[159][7] ;
 wire \cur_mb_mem[15][0] ;
 wire \cur_mb_mem[15][1] ;
 wire \cur_mb_mem[15][2] ;
 wire \cur_mb_mem[15][3] ;
 wire \cur_mb_mem[15][4] ;
 wire \cur_mb_mem[15][5] ;
 wire \cur_mb_mem[15][6] ;
 wire \cur_mb_mem[15][7] ;
 wire \cur_mb_mem[160][0] ;
 wire \cur_mb_mem[160][1] ;
 wire \cur_mb_mem[160][2] ;
 wire \cur_mb_mem[160][3] ;
 wire \cur_mb_mem[160][4] ;
 wire \cur_mb_mem[160][5] ;
 wire \cur_mb_mem[160][6] ;
 wire \cur_mb_mem[160][7] ;
 wire \cur_mb_mem[161][0] ;
 wire \cur_mb_mem[161][1] ;
 wire \cur_mb_mem[161][2] ;
 wire \cur_mb_mem[161][3] ;
 wire \cur_mb_mem[161][4] ;
 wire \cur_mb_mem[161][5] ;
 wire \cur_mb_mem[161][6] ;
 wire \cur_mb_mem[161][7] ;
 wire \cur_mb_mem[162][0] ;
 wire \cur_mb_mem[162][1] ;
 wire \cur_mb_mem[162][2] ;
 wire \cur_mb_mem[162][3] ;
 wire \cur_mb_mem[162][4] ;
 wire \cur_mb_mem[162][5] ;
 wire \cur_mb_mem[162][6] ;
 wire \cur_mb_mem[162][7] ;
 wire \cur_mb_mem[163][0] ;
 wire \cur_mb_mem[163][1] ;
 wire \cur_mb_mem[163][2] ;
 wire \cur_mb_mem[163][3] ;
 wire \cur_mb_mem[163][4] ;
 wire \cur_mb_mem[163][5] ;
 wire \cur_mb_mem[163][6] ;
 wire \cur_mb_mem[163][7] ;
 wire \cur_mb_mem[164][0] ;
 wire \cur_mb_mem[164][1] ;
 wire \cur_mb_mem[164][2] ;
 wire \cur_mb_mem[164][3] ;
 wire \cur_mb_mem[164][4] ;
 wire \cur_mb_mem[164][5] ;
 wire \cur_mb_mem[164][6] ;
 wire \cur_mb_mem[164][7] ;
 wire \cur_mb_mem[165][0] ;
 wire \cur_mb_mem[165][1] ;
 wire \cur_mb_mem[165][2] ;
 wire \cur_mb_mem[165][3] ;
 wire \cur_mb_mem[165][4] ;
 wire \cur_mb_mem[165][5] ;
 wire \cur_mb_mem[165][6] ;
 wire \cur_mb_mem[165][7] ;
 wire \cur_mb_mem[166][0] ;
 wire \cur_mb_mem[166][1] ;
 wire \cur_mb_mem[166][2] ;
 wire \cur_mb_mem[166][3] ;
 wire \cur_mb_mem[166][4] ;
 wire \cur_mb_mem[166][5] ;
 wire \cur_mb_mem[166][6] ;
 wire \cur_mb_mem[166][7] ;
 wire \cur_mb_mem[167][0] ;
 wire \cur_mb_mem[167][1] ;
 wire \cur_mb_mem[167][2] ;
 wire \cur_mb_mem[167][3] ;
 wire \cur_mb_mem[167][4] ;
 wire \cur_mb_mem[167][5] ;
 wire \cur_mb_mem[167][6] ;
 wire \cur_mb_mem[167][7] ;
 wire \cur_mb_mem[168][0] ;
 wire \cur_mb_mem[168][1] ;
 wire \cur_mb_mem[168][2] ;
 wire \cur_mb_mem[168][3] ;
 wire \cur_mb_mem[168][4] ;
 wire \cur_mb_mem[168][5] ;
 wire \cur_mb_mem[168][6] ;
 wire \cur_mb_mem[168][7] ;
 wire \cur_mb_mem[169][0] ;
 wire \cur_mb_mem[169][1] ;
 wire \cur_mb_mem[169][2] ;
 wire \cur_mb_mem[169][3] ;
 wire \cur_mb_mem[169][4] ;
 wire \cur_mb_mem[169][5] ;
 wire \cur_mb_mem[169][6] ;
 wire \cur_mb_mem[169][7] ;
 wire \cur_mb_mem[16][0] ;
 wire \cur_mb_mem[16][1] ;
 wire \cur_mb_mem[16][2] ;
 wire \cur_mb_mem[16][3] ;
 wire \cur_mb_mem[16][4] ;
 wire \cur_mb_mem[16][5] ;
 wire \cur_mb_mem[16][6] ;
 wire \cur_mb_mem[16][7] ;
 wire \cur_mb_mem[170][0] ;
 wire \cur_mb_mem[170][1] ;
 wire \cur_mb_mem[170][2] ;
 wire \cur_mb_mem[170][3] ;
 wire \cur_mb_mem[170][4] ;
 wire \cur_mb_mem[170][5] ;
 wire \cur_mb_mem[170][6] ;
 wire \cur_mb_mem[170][7] ;
 wire \cur_mb_mem[171][0] ;
 wire \cur_mb_mem[171][1] ;
 wire \cur_mb_mem[171][2] ;
 wire \cur_mb_mem[171][3] ;
 wire \cur_mb_mem[171][4] ;
 wire \cur_mb_mem[171][5] ;
 wire \cur_mb_mem[171][6] ;
 wire \cur_mb_mem[171][7] ;
 wire \cur_mb_mem[172][0] ;
 wire \cur_mb_mem[172][1] ;
 wire \cur_mb_mem[172][2] ;
 wire \cur_mb_mem[172][3] ;
 wire \cur_mb_mem[172][4] ;
 wire \cur_mb_mem[172][5] ;
 wire \cur_mb_mem[172][6] ;
 wire \cur_mb_mem[172][7] ;
 wire \cur_mb_mem[173][0] ;
 wire \cur_mb_mem[173][1] ;
 wire \cur_mb_mem[173][2] ;
 wire \cur_mb_mem[173][3] ;
 wire \cur_mb_mem[173][4] ;
 wire \cur_mb_mem[173][5] ;
 wire \cur_mb_mem[173][6] ;
 wire \cur_mb_mem[173][7] ;
 wire \cur_mb_mem[174][0] ;
 wire \cur_mb_mem[174][1] ;
 wire \cur_mb_mem[174][2] ;
 wire \cur_mb_mem[174][3] ;
 wire \cur_mb_mem[174][4] ;
 wire \cur_mb_mem[174][5] ;
 wire \cur_mb_mem[174][6] ;
 wire \cur_mb_mem[174][7] ;
 wire \cur_mb_mem[175][0] ;
 wire \cur_mb_mem[175][1] ;
 wire \cur_mb_mem[175][2] ;
 wire \cur_mb_mem[175][3] ;
 wire \cur_mb_mem[175][4] ;
 wire \cur_mb_mem[175][5] ;
 wire \cur_mb_mem[175][6] ;
 wire \cur_mb_mem[175][7] ;
 wire \cur_mb_mem[176][0] ;
 wire \cur_mb_mem[176][1] ;
 wire \cur_mb_mem[176][2] ;
 wire \cur_mb_mem[176][3] ;
 wire \cur_mb_mem[176][4] ;
 wire \cur_mb_mem[176][5] ;
 wire \cur_mb_mem[176][6] ;
 wire \cur_mb_mem[176][7] ;
 wire \cur_mb_mem[177][0] ;
 wire \cur_mb_mem[177][1] ;
 wire \cur_mb_mem[177][2] ;
 wire \cur_mb_mem[177][3] ;
 wire \cur_mb_mem[177][4] ;
 wire \cur_mb_mem[177][5] ;
 wire \cur_mb_mem[177][6] ;
 wire \cur_mb_mem[177][7] ;
 wire \cur_mb_mem[178][0] ;
 wire \cur_mb_mem[178][1] ;
 wire \cur_mb_mem[178][2] ;
 wire \cur_mb_mem[178][3] ;
 wire \cur_mb_mem[178][4] ;
 wire \cur_mb_mem[178][5] ;
 wire \cur_mb_mem[178][6] ;
 wire \cur_mb_mem[178][7] ;
 wire \cur_mb_mem[179][0] ;
 wire \cur_mb_mem[179][1] ;
 wire \cur_mb_mem[179][2] ;
 wire \cur_mb_mem[179][3] ;
 wire \cur_mb_mem[179][4] ;
 wire \cur_mb_mem[179][5] ;
 wire \cur_mb_mem[179][6] ;
 wire \cur_mb_mem[179][7] ;
 wire \cur_mb_mem[17][0] ;
 wire \cur_mb_mem[17][1] ;
 wire \cur_mb_mem[17][2] ;
 wire \cur_mb_mem[17][3] ;
 wire \cur_mb_mem[17][4] ;
 wire \cur_mb_mem[17][5] ;
 wire \cur_mb_mem[17][6] ;
 wire \cur_mb_mem[17][7] ;
 wire \cur_mb_mem[180][0] ;
 wire \cur_mb_mem[180][1] ;
 wire \cur_mb_mem[180][2] ;
 wire \cur_mb_mem[180][3] ;
 wire \cur_mb_mem[180][4] ;
 wire \cur_mb_mem[180][5] ;
 wire \cur_mb_mem[180][6] ;
 wire \cur_mb_mem[180][7] ;
 wire \cur_mb_mem[181][0] ;
 wire \cur_mb_mem[181][1] ;
 wire \cur_mb_mem[181][2] ;
 wire \cur_mb_mem[181][3] ;
 wire \cur_mb_mem[181][4] ;
 wire \cur_mb_mem[181][5] ;
 wire \cur_mb_mem[181][6] ;
 wire \cur_mb_mem[181][7] ;
 wire \cur_mb_mem[182][0] ;
 wire \cur_mb_mem[182][1] ;
 wire \cur_mb_mem[182][2] ;
 wire \cur_mb_mem[182][3] ;
 wire \cur_mb_mem[182][4] ;
 wire \cur_mb_mem[182][5] ;
 wire \cur_mb_mem[182][6] ;
 wire \cur_mb_mem[182][7] ;
 wire \cur_mb_mem[183][0] ;
 wire \cur_mb_mem[183][1] ;
 wire \cur_mb_mem[183][2] ;
 wire \cur_mb_mem[183][3] ;
 wire \cur_mb_mem[183][4] ;
 wire \cur_mb_mem[183][5] ;
 wire \cur_mb_mem[183][6] ;
 wire \cur_mb_mem[183][7] ;
 wire \cur_mb_mem[184][0] ;
 wire \cur_mb_mem[184][1] ;
 wire \cur_mb_mem[184][2] ;
 wire \cur_mb_mem[184][3] ;
 wire \cur_mb_mem[184][4] ;
 wire \cur_mb_mem[184][5] ;
 wire \cur_mb_mem[184][6] ;
 wire \cur_mb_mem[184][7] ;
 wire \cur_mb_mem[185][0] ;
 wire \cur_mb_mem[185][1] ;
 wire \cur_mb_mem[185][2] ;
 wire \cur_mb_mem[185][3] ;
 wire \cur_mb_mem[185][4] ;
 wire \cur_mb_mem[185][5] ;
 wire \cur_mb_mem[185][6] ;
 wire \cur_mb_mem[185][7] ;
 wire \cur_mb_mem[186][0] ;
 wire \cur_mb_mem[186][1] ;
 wire \cur_mb_mem[186][2] ;
 wire \cur_mb_mem[186][3] ;
 wire \cur_mb_mem[186][4] ;
 wire \cur_mb_mem[186][5] ;
 wire \cur_mb_mem[186][6] ;
 wire \cur_mb_mem[186][7] ;
 wire \cur_mb_mem[187][0] ;
 wire \cur_mb_mem[187][1] ;
 wire \cur_mb_mem[187][2] ;
 wire \cur_mb_mem[187][3] ;
 wire \cur_mb_mem[187][4] ;
 wire \cur_mb_mem[187][5] ;
 wire \cur_mb_mem[187][6] ;
 wire \cur_mb_mem[187][7] ;
 wire \cur_mb_mem[188][0] ;
 wire \cur_mb_mem[188][1] ;
 wire \cur_mb_mem[188][2] ;
 wire \cur_mb_mem[188][3] ;
 wire \cur_mb_mem[188][4] ;
 wire \cur_mb_mem[188][5] ;
 wire \cur_mb_mem[188][6] ;
 wire \cur_mb_mem[188][7] ;
 wire \cur_mb_mem[189][0] ;
 wire \cur_mb_mem[189][1] ;
 wire \cur_mb_mem[189][2] ;
 wire \cur_mb_mem[189][3] ;
 wire \cur_mb_mem[189][4] ;
 wire \cur_mb_mem[189][5] ;
 wire \cur_mb_mem[189][6] ;
 wire \cur_mb_mem[189][7] ;
 wire \cur_mb_mem[18][0] ;
 wire \cur_mb_mem[18][1] ;
 wire \cur_mb_mem[18][2] ;
 wire \cur_mb_mem[18][3] ;
 wire \cur_mb_mem[18][4] ;
 wire \cur_mb_mem[18][5] ;
 wire \cur_mb_mem[18][6] ;
 wire \cur_mb_mem[18][7] ;
 wire \cur_mb_mem[190][0] ;
 wire \cur_mb_mem[190][1] ;
 wire \cur_mb_mem[190][2] ;
 wire \cur_mb_mem[190][3] ;
 wire \cur_mb_mem[190][4] ;
 wire \cur_mb_mem[190][5] ;
 wire \cur_mb_mem[190][6] ;
 wire \cur_mb_mem[190][7] ;
 wire \cur_mb_mem[191][0] ;
 wire \cur_mb_mem[191][1] ;
 wire \cur_mb_mem[191][2] ;
 wire \cur_mb_mem[191][3] ;
 wire \cur_mb_mem[191][4] ;
 wire \cur_mb_mem[191][5] ;
 wire \cur_mb_mem[191][6] ;
 wire \cur_mb_mem[191][7] ;
 wire \cur_mb_mem[192][0] ;
 wire \cur_mb_mem[192][1] ;
 wire \cur_mb_mem[192][2] ;
 wire \cur_mb_mem[192][3] ;
 wire \cur_mb_mem[192][4] ;
 wire \cur_mb_mem[192][5] ;
 wire \cur_mb_mem[192][6] ;
 wire \cur_mb_mem[192][7] ;
 wire \cur_mb_mem[193][0] ;
 wire \cur_mb_mem[193][1] ;
 wire \cur_mb_mem[193][2] ;
 wire \cur_mb_mem[193][3] ;
 wire \cur_mb_mem[193][4] ;
 wire \cur_mb_mem[193][5] ;
 wire \cur_mb_mem[193][6] ;
 wire \cur_mb_mem[193][7] ;
 wire \cur_mb_mem[194][0] ;
 wire \cur_mb_mem[194][1] ;
 wire \cur_mb_mem[194][2] ;
 wire \cur_mb_mem[194][3] ;
 wire \cur_mb_mem[194][4] ;
 wire \cur_mb_mem[194][5] ;
 wire \cur_mb_mem[194][6] ;
 wire \cur_mb_mem[194][7] ;
 wire \cur_mb_mem[195][0] ;
 wire \cur_mb_mem[195][1] ;
 wire \cur_mb_mem[195][2] ;
 wire \cur_mb_mem[195][3] ;
 wire \cur_mb_mem[195][4] ;
 wire \cur_mb_mem[195][5] ;
 wire \cur_mb_mem[195][6] ;
 wire \cur_mb_mem[195][7] ;
 wire \cur_mb_mem[196][0] ;
 wire \cur_mb_mem[196][1] ;
 wire \cur_mb_mem[196][2] ;
 wire \cur_mb_mem[196][3] ;
 wire \cur_mb_mem[196][4] ;
 wire \cur_mb_mem[196][5] ;
 wire \cur_mb_mem[196][6] ;
 wire \cur_mb_mem[196][7] ;
 wire \cur_mb_mem[197][0] ;
 wire \cur_mb_mem[197][1] ;
 wire \cur_mb_mem[197][2] ;
 wire \cur_mb_mem[197][3] ;
 wire \cur_mb_mem[197][4] ;
 wire \cur_mb_mem[197][5] ;
 wire \cur_mb_mem[197][6] ;
 wire \cur_mb_mem[197][7] ;
 wire \cur_mb_mem[198][0] ;
 wire \cur_mb_mem[198][1] ;
 wire \cur_mb_mem[198][2] ;
 wire \cur_mb_mem[198][3] ;
 wire \cur_mb_mem[198][4] ;
 wire \cur_mb_mem[198][5] ;
 wire \cur_mb_mem[198][6] ;
 wire \cur_mb_mem[198][7] ;
 wire \cur_mb_mem[199][0] ;
 wire \cur_mb_mem[199][1] ;
 wire \cur_mb_mem[199][2] ;
 wire \cur_mb_mem[199][3] ;
 wire \cur_mb_mem[199][4] ;
 wire \cur_mb_mem[199][5] ;
 wire \cur_mb_mem[199][6] ;
 wire \cur_mb_mem[199][7] ;
 wire \cur_mb_mem[19][0] ;
 wire \cur_mb_mem[19][1] ;
 wire \cur_mb_mem[19][2] ;
 wire \cur_mb_mem[19][3] ;
 wire \cur_mb_mem[19][4] ;
 wire \cur_mb_mem[19][5] ;
 wire \cur_mb_mem[19][6] ;
 wire \cur_mb_mem[19][7] ;
 wire \cur_mb_mem[1][0] ;
 wire \cur_mb_mem[1][1] ;
 wire \cur_mb_mem[1][2] ;
 wire \cur_mb_mem[1][3] ;
 wire \cur_mb_mem[1][4] ;
 wire \cur_mb_mem[1][5] ;
 wire \cur_mb_mem[1][6] ;
 wire \cur_mb_mem[1][7] ;
 wire \cur_mb_mem[200][0] ;
 wire \cur_mb_mem[200][1] ;
 wire \cur_mb_mem[200][2] ;
 wire \cur_mb_mem[200][3] ;
 wire \cur_mb_mem[200][4] ;
 wire \cur_mb_mem[200][5] ;
 wire \cur_mb_mem[200][6] ;
 wire \cur_mb_mem[200][7] ;
 wire \cur_mb_mem[201][0] ;
 wire \cur_mb_mem[201][1] ;
 wire \cur_mb_mem[201][2] ;
 wire \cur_mb_mem[201][3] ;
 wire \cur_mb_mem[201][4] ;
 wire \cur_mb_mem[201][5] ;
 wire \cur_mb_mem[201][6] ;
 wire \cur_mb_mem[201][7] ;
 wire \cur_mb_mem[202][0] ;
 wire \cur_mb_mem[202][1] ;
 wire \cur_mb_mem[202][2] ;
 wire \cur_mb_mem[202][3] ;
 wire \cur_mb_mem[202][4] ;
 wire \cur_mb_mem[202][5] ;
 wire \cur_mb_mem[202][6] ;
 wire \cur_mb_mem[202][7] ;
 wire \cur_mb_mem[203][0] ;
 wire \cur_mb_mem[203][1] ;
 wire \cur_mb_mem[203][2] ;
 wire \cur_mb_mem[203][3] ;
 wire \cur_mb_mem[203][4] ;
 wire \cur_mb_mem[203][5] ;
 wire \cur_mb_mem[203][6] ;
 wire \cur_mb_mem[203][7] ;
 wire \cur_mb_mem[204][0] ;
 wire \cur_mb_mem[204][1] ;
 wire \cur_mb_mem[204][2] ;
 wire \cur_mb_mem[204][3] ;
 wire \cur_mb_mem[204][4] ;
 wire \cur_mb_mem[204][5] ;
 wire \cur_mb_mem[204][6] ;
 wire \cur_mb_mem[204][7] ;
 wire \cur_mb_mem[205][0] ;
 wire \cur_mb_mem[205][1] ;
 wire \cur_mb_mem[205][2] ;
 wire \cur_mb_mem[205][3] ;
 wire \cur_mb_mem[205][4] ;
 wire \cur_mb_mem[205][5] ;
 wire \cur_mb_mem[205][6] ;
 wire \cur_mb_mem[205][7] ;
 wire \cur_mb_mem[206][0] ;
 wire \cur_mb_mem[206][1] ;
 wire \cur_mb_mem[206][2] ;
 wire \cur_mb_mem[206][3] ;
 wire \cur_mb_mem[206][4] ;
 wire \cur_mb_mem[206][5] ;
 wire \cur_mb_mem[206][6] ;
 wire \cur_mb_mem[206][7] ;
 wire \cur_mb_mem[207][0] ;
 wire \cur_mb_mem[207][1] ;
 wire \cur_mb_mem[207][2] ;
 wire \cur_mb_mem[207][3] ;
 wire \cur_mb_mem[207][4] ;
 wire \cur_mb_mem[207][5] ;
 wire \cur_mb_mem[207][6] ;
 wire \cur_mb_mem[207][7] ;
 wire \cur_mb_mem[208][0] ;
 wire \cur_mb_mem[208][1] ;
 wire \cur_mb_mem[208][2] ;
 wire \cur_mb_mem[208][3] ;
 wire \cur_mb_mem[208][4] ;
 wire \cur_mb_mem[208][5] ;
 wire \cur_mb_mem[208][6] ;
 wire \cur_mb_mem[208][7] ;
 wire \cur_mb_mem[209][0] ;
 wire \cur_mb_mem[209][1] ;
 wire \cur_mb_mem[209][2] ;
 wire \cur_mb_mem[209][3] ;
 wire \cur_mb_mem[209][4] ;
 wire \cur_mb_mem[209][5] ;
 wire \cur_mb_mem[209][6] ;
 wire \cur_mb_mem[209][7] ;
 wire \cur_mb_mem[20][0] ;
 wire \cur_mb_mem[20][1] ;
 wire \cur_mb_mem[20][2] ;
 wire \cur_mb_mem[20][3] ;
 wire \cur_mb_mem[20][4] ;
 wire \cur_mb_mem[20][5] ;
 wire \cur_mb_mem[20][6] ;
 wire \cur_mb_mem[20][7] ;
 wire \cur_mb_mem[210][0] ;
 wire \cur_mb_mem[210][1] ;
 wire \cur_mb_mem[210][2] ;
 wire \cur_mb_mem[210][3] ;
 wire \cur_mb_mem[210][4] ;
 wire \cur_mb_mem[210][5] ;
 wire \cur_mb_mem[210][6] ;
 wire \cur_mb_mem[210][7] ;
 wire \cur_mb_mem[211][0] ;
 wire \cur_mb_mem[211][1] ;
 wire \cur_mb_mem[211][2] ;
 wire \cur_mb_mem[211][3] ;
 wire \cur_mb_mem[211][4] ;
 wire \cur_mb_mem[211][5] ;
 wire \cur_mb_mem[211][6] ;
 wire \cur_mb_mem[211][7] ;
 wire \cur_mb_mem[212][0] ;
 wire \cur_mb_mem[212][1] ;
 wire \cur_mb_mem[212][2] ;
 wire \cur_mb_mem[212][3] ;
 wire \cur_mb_mem[212][4] ;
 wire \cur_mb_mem[212][5] ;
 wire \cur_mb_mem[212][6] ;
 wire \cur_mb_mem[212][7] ;
 wire \cur_mb_mem[213][0] ;
 wire \cur_mb_mem[213][1] ;
 wire \cur_mb_mem[213][2] ;
 wire \cur_mb_mem[213][3] ;
 wire \cur_mb_mem[213][4] ;
 wire \cur_mb_mem[213][5] ;
 wire \cur_mb_mem[213][6] ;
 wire \cur_mb_mem[213][7] ;
 wire \cur_mb_mem[214][0] ;
 wire \cur_mb_mem[214][1] ;
 wire \cur_mb_mem[214][2] ;
 wire \cur_mb_mem[214][3] ;
 wire \cur_mb_mem[214][4] ;
 wire \cur_mb_mem[214][5] ;
 wire \cur_mb_mem[214][6] ;
 wire \cur_mb_mem[214][7] ;
 wire \cur_mb_mem[215][0] ;
 wire \cur_mb_mem[215][1] ;
 wire \cur_mb_mem[215][2] ;
 wire \cur_mb_mem[215][3] ;
 wire \cur_mb_mem[215][4] ;
 wire \cur_mb_mem[215][5] ;
 wire \cur_mb_mem[215][6] ;
 wire \cur_mb_mem[215][7] ;
 wire \cur_mb_mem[216][0] ;
 wire \cur_mb_mem[216][1] ;
 wire \cur_mb_mem[216][2] ;
 wire \cur_mb_mem[216][3] ;
 wire \cur_mb_mem[216][4] ;
 wire \cur_mb_mem[216][5] ;
 wire \cur_mb_mem[216][6] ;
 wire \cur_mb_mem[216][7] ;
 wire \cur_mb_mem[217][0] ;
 wire \cur_mb_mem[217][1] ;
 wire \cur_mb_mem[217][2] ;
 wire \cur_mb_mem[217][3] ;
 wire \cur_mb_mem[217][4] ;
 wire \cur_mb_mem[217][5] ;
 wire \cur_mb_mem[217][6] ;
 wire \cur_mb_mem[217][7] ;
 wire \cur_mb_mem[218][0] ;
 wire \cur_mb_mem[218][1] ;
 wire \cur_mb_mem[218][2] ;
 wire \cur_mb_mem[218][3] ;
 wire \cur_mb_mem[218][4] ;
 wire \cur_mb_mem[218][5] ;
 wire \cur_mb_mem[218][6] ;
 wire \cur_mb_mem[218][7] ;
 wire \cur_mb_mem[219][0] ;
 wire \cur_mb_mem[219][1] ;
 wire \cur_mb_mem[219][2] ;
 wire \cur_mb_mem[219][3] ;
 wire \cur_mb_mem[219][4] ;
 wire \cur_mb_mem[219][5] ;
 wire \cur_mb_mem[219][6] ;
 wire \cur_mb_mem[219][7] ;
 wire \cur_mb_mem[21][0] ;
 wire \cur_mb_mem[21][1] ;
 wire \cur_mb_mem[21][2] ;
 wire \cur_mb_mem[21][3] ;
 wire \cur_mb_mem[21][4] ;
 wire \cur_mb_mem[21][5] ;
 wire \cur_mb_mem[21][6] ;
 wire \cur_mb_mem[21][7] ;
 wire \cur_mb_mem[220][0] ;
 wire \cur_mb_mem[220][1] ;
 wire \cur_mb_mem[220][2] ;
 wire \cur_mb_mem[220][3] ;
 wire \cur_mb_mem[220][4] ;
 wire \cur_mb_mem[220][5] ;
 wire \cur_mb_mem[220][6] ;
 wire \cur_mb_mem[220][7] ;
 wire \cur_mb_mem[221][0] ;
 wire \cur_mb_mem[221][1] ;
 wire \cur_mb_mem[221][2] ;
 wire \cur_mb_mem[221][3] ;
 wire \cur_mb_mem[221][4] ;
 wire \cur_mb_mem[221][5] ;
 wire \cur_mb_mem[221][6] ;
 wire \cur_mb_mem[221][7] ;
 wire \cur_mb_mem[222][0] ;
 wire \cur_mb_mem[222][1] ;
 wire \cur_mb_mem[222][2] ;
 wire \cur_mb_mem[222][3] ;
 wire \cur_mb_mem[222][4] ;
 wire \cur_mb_mem[222][5] ;
 wire \cur_mb_mem[222][6] ;
 wire \cur_mb_mem[222][7] ;
 wire \cur_mb_mem[223][0] ;
 wire \cur_mb_mem[223][1] ;
 wire \cur_mb_mem[223][2] ;
 wire \cur_mb_mem[223][3] ;
 wire \cur_mb_mem[223][4] ;
 wire \cur_mb_mem[223][5] ;
 wire \cur_mb_mem[223][6] ;
 wire \cur_mb_mem[223][7] ;
 wire \cur_mb_mem[224][0] ;
 wire \cur_mb_mem[224][1] ;
 wire \cur_mb_mem[224][2] ;
 wire \cur_mb_mem[224][3] ;
 wire \cur_mb_mem[224][4] ;
 wire \cur_mb_mem[224][5] ;
 wire \cur_mb_mem[224][6] ;
 wire \cur_mb_mem[224][7] ;
 wire \cur_mb_mem[225][0] ;
 wire \cur_mb_mem[225][1] ;
 wire \cur_mb_mem[225][2] ;
 wire \cur_mb_mem[225][3] ;
 wire \cur_mb_mem[225][4] ;
 wire \cur_mb_mem[225][5] ;
 wire \cur_mb_mem[225][6] ;
 wire \cur_mb_mem[225][7] ;
 wire \cur_mb_mem[226][0] ;
 wire \cur_mb_mem[226][1] ;
 wire \cur_mb_mem[226][2] ;
 wire \cur_mb_mem[226][3] ;
 wire \cur_mb_mem[226][4] ;
 wire \cur_mb_mem[226][5] ;
 wire \cur_mb_mem[226][6] ;
 wire \cur_mb_mem[226][7] ;
 wire \cur_mb_mem[227][0] ;
 wire \cur_mb_mem[227][1] ;
 wire \cur_mb_mem[227][2] ;
 wire \cur_mb_mem[227][3] ;
 wire \cur_mb_mem[227][4] ;
 wire \cur_mb_mem[227][5] ;
 wire \cur_mb_mem[227][6] ;
 wire \cur_mb_mem[227][7] ;
 wire \cur_mb_mem[228][0] ;
 wire \cur_mb_mem[228][1] ;
 wire \cur_mb_mem[228][2] ;
 wire \cur_mb_mem[228][3] ;
 wire \cur_mb_mem[228][4] ;
 wire \cur_mb_mem[228][5] ;
 wire \cur_mb_mem[228][6] ;
 wire \cur_mb_mem[228][7] ;
 wire \cur_mb_mem[229][0] ;
 wire \cur_mb_mem[229][1] ;
 wire \cur_mb_mem[229][2] ;
 wire \cur_mb_mem[229][3] ;
 wire \cur_mb_mem[229][4] ;
 wire \cur_mb_mem[229][5] ;
 wire \cur_mb_mem[229][6] ;
 wire \cur_mb_mem[229][7] ;
 wire \cur_mb_mem[22][0] ;
 wire \cur_mb_mem[22][1] ;
 wire \cur_mb_mem[22][2] ;
 wire \cur_mb_mem[22][3] ;
 wire \cur_mb_mem[22][4] ;
 wire \cur_mb_mem[22][5] ;
 wire \cur_mb_mem[22][6] ;
 wire \cur_mb_mem[22][7] ;
 wire \cur_mb_mem[230][0] ;
 wire \cur_mb_mem[230][1] ;
 wire \cur_mb_mem[230][2] ;
 wire \cur_mb_mem[230][3] ;
 wire \cur_mb_mem[230][4] ;
 wire \cur_mb_mem[230][5] ;
 wire \cur_mb_mem[230][6] ;
 wire \cur_mb_mem[230][7] ;
 wire \cur_mb_mem[231][0] ;
 wire \cur_mb_mem[231][1] ;
 wire \cur_mb_mem[231][2] ;
 wire \cur_mb_mem[231][3] ;
 wire \cur_mb_mem[231][4] ;
 wire \cur_mb_mem[231][5] ;
 wire \cur_mb_mem[231][6] ;
 wire \cur_mb_mem[231][7] ;
 wire \cur_mb_mem[232][0] ;
 wire \cur_mb_mem[232][1] ;
 wire \cur_mb_mem[232][2] ;
 wire \cur_mb_mem[232][3] ;
 wire \cur_mb_mem[232][4] ;
 wire \cur_mb_mem[232][5] ;
 wire \cur_mb_mem[232][6] ;
 wire \cur_mb_mem[232][7] ;
 wire \cur_mb_mem[233][0] ;
 wire \cur_mb_mem[233][1] ;
 wire \cur_mb_mem[233][2] ;
 wire \cur_mb_mem[233][3] ;
 wire \cur_mb_mem[233][4] ;
 wire \cur_mb_mem[233][5] ;
 wire \cur_mb_mem[233][6] ;
 wire \cur_mb_mem[233][7] ;
 wire \cur_mb_mem[234][0] ;
 wire \cur_mb_mem[234][1] ;
 wire \cur_mb_mem[234][2] ;
 wire \cur_mb_mem[234][3] ;
 wire \cur_mb_mem[234][4] ;
 wire \cur_mb_mem[234][5] ;
 wire \cur_mb_mem[234][6] ;
 wire \cur_mb_mem[234][7] ;
 wire \cur_mb_mem[235][0] ;
 wire \cur_mb_mem[235][1] ;
 wire \cur_mb_mem[235][2] ;
 wire \cur_mb_mem[235][3] ;
 wire \cur_mb_mem[235][4] ;
 wire \cur_mb_mem[235][5] ;
 wire \cur_mb_mem[235][6] ;
 wire \cur_mb_mem[235][7] ;
 wire \cur_mb_mem[236][0] ;
 wire \cur_mb_mem[236][1] ;
 wire \cur_mb_mem[236][2] ;
 wire \cur_mb_mem[236][3] ;
 wire \cur_mb_mem[236][4] ;
 wire \cur_mb_mem[236][5] ;
 wire \cur_mb_mem[236][6] ;
 wire \cur_mb_mem[236][7] ;
 wire \cur_mb_mem[237][0] ;
 wire \cur_mb_mem[237][1] ;
 wire \cur_mb_mem[237][2] ;
 wire \cur_mb_mem[237][3] ;
 wire \cur_mb_mem[237][4] ;
 wire \cur_mb_mem[237][5] ;
 wire \cur_mb_mem[237][6] ;
 wire \cur_mb_mem[237][7] ;
 wire \cur_mb_mem[238][0] ;
 wire \cur_mb_mem[238][1] ;
 wire \cur_mb_mem[238][2] ;
 wire \cur_mb_mem[238][3] ;
 wire \cur_mb_mem[238][4] ;
 wire \cur_mb_mem[238][5] ;
 wire \cur_mb_mem[238][6] ;
 wire \cur_mb_mem[238][7] ;
 wire \cur_mb_mem[239][0] ;
 wire \cur_mb_mem[239][1] ;
 wire \cur_mb_mem[239][2] ;
 wire \cur_mb_mem[239][3] ;
 wire \cur_mb_mem[239][4] ;
 wire \cur_mb_mem[239][5] ;
 wire \cur_mb_mem[239][6] ;
 wire \cur_mb_mem[239][7] ;
 wire \cur_mb_mem[23][0] ;
 wire \cur_mb_mem[23][1] ;
 wire \cur_mb_mem[23][2] ;
 wire \cur_mb_mem[23][3] ;
 wire \cur_mb_mem[23][4] ;
 wire \cur_mb_mem[23][5] ;
 wire \cur_mb_mem[23][6] ;
 wire \cur_mb_mem[23][7] ;
 wire \cur_mb_mem[240][0] ;
 wire \cur_mb_mem[240][1] ;
 wire \cur_mb_mem[240][2] ;
 wire \cur_mb_mem[240][3] ;
 wire \cur_mb_mem[240][4] ;
 wire \cur_mb_mem[240][5] ;
 wire \cur_mb_mem[240][6] ;
 wire \cur_mb_mem[240][7] ;
 wire \cur_mb_mem[241][0] ;
 wire \cur_mb_mem[241][1] ;
 wire \cur_mb_mem[241][2] ;
 wire \cur_mb_mem[241][3] ;
 wire \cur_mb_mem[241][4] ;
 wire \cur_mb_mem[241][5] ;
 wire \cur_mb_mem[241][6] ;
 wire \cur_mb_mem[241][7] ;
 wire \cur_mb_mem[242][0] ;
 wire \cur_mb_mem[242][1] ;
 wire \cur_mb_mem[242][2] ;
 wire \cur_mb_mem[242][3] ;
 wire \cur_mb_mem[242][4] ;
 wire \cur_mb_mem[242][5] ;
 wire \cur_mb_mem[242][6] ;
 wire \cur_mb_mem[242][7] ;
 wire \cur_mb_mem[243][0] ;
 wire \cur_mb_mem[243][1] ;
 wire \cur_mb_mem[243][2] ;
 wire \cur_mb_mem[243][3] ;
 wire \cur_mb_mem[243][4] ;
 wire \cur_mb_mem[243][5] ;
 wire \cur_mb_mem[243][6] ;
 wire \cur_mb_mem[243][7] ;
 wire \cur_mb_mem[244][0] ;
 wire \cur_mb_mem[244][1] ;
 wire \cur_mb_mem[244][2] ;
 wire \cur_mb_mem[244][3] ;
 wire \cur_mb_mem[244][4] ;
 wire \cur_mb_mem[244][5] ;
 wire \cur_mb_mem[244][6] ;
 wire \cur_mb_mem[244][7] ;
 wire \cur_mb_mem[245][0] ;
 wire \cur_mb_mem[245][1] ;
 wire \cur_mb_mem[245][2] ;
 wire \cur_mb_mem[245][3] ;
 wire \cur_mb_mem[245][4] ;
 wire \cur_mb_mem[245][5] ;
 wire \cur_mb_mem[245][6] ;
 wire \cur_mb_mem[245][7] ;
 wire \cur_mb_mem[246][0] ;
 wire \cur_mb_mem[246][1] ;
 wire \cur_mb_mem[246][2] ;
 wire \cur_mb_mem[246][3] ;
 wire \cur_mb_mem[246][4] ;
 wire \cur_mb_mem[246][5] ;
 wire \cur_mb_mem[246][6] ;
 wire \cur_mb_mem[246][7] ;
 wire \cur_mb_mem[247][0] ;
 wire \cur_mb_mem[247][1] ;
 wire \cur_mb_mem[247][2] ;
 wire \cur_mb_mem[247][3] ;
 wire \cur_mb_mem[247][4] ;
 wire \cur_mb_mem[247][5] ;
 wire \cur_mb_mem[247][6] ;
 wire \cur_mb_mem[247][7] ;
 wire \cur_mb_mem[248][0] ;
 wire \cur_mb_mem[248][1] ;
 wire \cur_mb_mem[248][2] ;
 wire \cur_mb_mem[248][3] ;
 wire \cur_mb_mem[248][4] ;
 wire \cur_mb_mem[248][5] ;
 wire \cur_mb_mem[248][6] ;
 wire \cur_mb_mem[248][7] ;
 wire \cur_mb_mem[249][0] ;
 wire \cur_mb_mem[249][1] ;
 wire \cur_mb_mem[249][2] ;
 wire \cur_mb_mem[249][3] ;
 wire \cur_mb_mem[249][4] ;
 wire \cur_mb_mem[249][5] ;
 wire \cur_mb_mem[249][6] ;
 wire \cur_mb_mem[249][7] ;
 wire \cur_mb_mem[24][0] ;
 wire \cur_mb_mem[24][1] ;
 wire \cur_mb_mem[24][2] ;
 wire \cur_mb_mem[24][3] ;
 wire \cur_mb_mem[24][4] ;
 wire \cur_mb_mem[24][5] ;
 wire \cur_mb_mem[24][6] ;
 wire \cur_mb_mem[24][7] ;
 wire \cur_mb_mem[250][0] ;
 wire \cur_mb_mem[250][1] ;
 wire \cur_mb_mem[250][2] ;
 wire \cur_mb_mem[250][3] ;
 wire \cur_mb_mem[250][4] ;
 wire \cur_mb_mem[250][5] ;
 wire \cur_mb_mem[250][6] ;
 wire \cur_mb_mem[250][7] ;
 wire \cur_mb_mem[251][0] ;
 wire \cur_mb_mem[251][1] ;
 wire \cur_mb_mem[251][2] ;
 wire \cur_mb_mem[251][3] ;
 wire \cur_mb_mem[251][4] ;
 wire \cur_mb_mem[251][5] ;
 wire \cur_mb_mem[251][6] ;
 wire \cur_mb_mem[251][7] ;
 wire \cur_mb_mem[252][0] ;
 wire \cur_mb_mem[252][1] ;
 wire \cur_mb_mem[252][2] ;
 wire \cur_mb_mem[252][3] ;
 wire \cur_mb_mem[252][4] ;
 wire \cur_mb_mem[252][5] ;
 wire \cur_mb_mem[252][6] ;
 wire \cur_mb_mem[252][7] ;
 wire \cur_mb_mem[253][0] ;
 wire \cur_mb_mem[253][1] ;
 wire \cur_mb_mem[253][2] ;
 wire \cur_mb_mem[253][3] ;
 wire \cur_mb_mem[253][4] ;
 wire \cur_mb_mem[253][5] ;
 wire \cur_mb_mem[253][6] ;
 wire \cur_mb_mem[253][7] ;
 wire \cur_mb_mem[254][0] ;
 wire \cur_mb_mem[254][1] ;
 wire \cur_mb_mem[254][2] ;
 wire \cur_mb_mem[254][3] ;
 wire \cur_mb_mem[254][4] ;
 wire \cur_mb_mem[254][5] ;
 wire \cur_mb_mem[254][6] ;
 wire \cur_mb_mem[254][7] ;
 wire \cur_mb_mem[255][0] ;
 wire \cur_mb_mem[255][1] ;
 wire \cur_mb_mem[255][2] ;
 wire \cur_mb_mem[255][3] ;
 wire \cur_mb_mem[255][4] ;
 wire \cur_mb_mem[255][5] ;
 wire \cur_mb_mem[255][6] ;
 wire \cur_mb_mem[255][7] ;
 wire \cur_mb_mem[25][0] ;
 wire \cur_mb_mem[25][1] ;
 wire \cur_mb_mem[25][2] ;
 wire \cur_mb_mem[25][3] ;
 wire \cur_mb_mem[25][4] ;
 wire \cur_mb_mem[25][5] ;
 wire \cur_mb_mem[25][6] ;
 wire \cur_mb_mem[25][7] ;
 wire \cur_mb_mem[26][0] ;
 wire \cur_mb_mem[26][1] ;
 wire \cur_mb_mem[26][2] ;
 wire \cur_mb_mem[26][3] ;
 wire \cur_mb_mem[26][4] ;
 wire \cur_mb_mem[26][5] ;
 wire \cur_mb_mem[26][6] ;
 wire \cur_mb_mem[26][7] ;
 wire \cur_mb_mem[27][0] ;
 wire \cur_mb_mem[27][1] ;
 wire \cur_mb_mem[27][2] ;
 wire \cur_mb_mem[27][3] ;
 wire \cur_mb_mem[27][4] ;
 wire \cur_mb_mem[27][5] ;
 wire \cur_mb_mem[27][6] ;
 wire \cur_mb_mem[27][7] ;
 wire \cur_mb_mem[28][0] ;
 wire \cur_mb_mem[28][1] ;
 wire \cur_mb_mem[28][2] ;
 wire \cur_mb_mem[28][3] ;
 wire \cur_mb_mem[28][4] ;
 wire \cur_mb_mem[28][5] ;
 wire \cur_mb_mem[28][6] ;
 wire \cur_mb_mem[28][7] ;
 wire \cur_mb_mem[29][0] ;
 wire \cur_mb_mem[29][1] ;
 wire \cur_mb_mem[29][2] ;
 wire \cur_mb_mem[29][3] ;
 wire \cur_mb_mem[29][4] ;
 wire \cur_mb_mem[29][5] ;
 wire \cur_mb_mem[29][6] ;
 wire \cur_mb_mem[29][7] ;
 wire \cur_mb_mem[2][0] ;
 wire \cur_mb_mem[2][1] ;
 wire \cur_mb_mem[2][2] ;
 wire \cur_mb_mem[2][3] ;
 wire \cur_mb_mem[2][4] ;
 wire \cur_mb_mem[2][5] ;
 wire \cur_mb_mem[2][6] ;
 wire \cur_mb_mem[2][7] ;
 wire \cur_mb_mem[30][0] ;
 wire \cur_mb_mem[30][1] ;
 wire \cur_mb_mem[30][2] ;
 wire \cur_mb_mem[30][3] ;
 wire \cur_mb_mem[30][4] ;
 wire \cur_mb_mem[30][5] ;
 wire \cur_mb_mem[30][6] ;
 wire \cur_mb_mem[30][7] ;
 wire \cur_mb_mem[31][0] ;
 wire \cur_mb_mem[31][1] ;
 wire \cur_mb_mem[31][2] ;
 wire \cur_mb_mem[31][3] ;
 wire \cur_mb_mem[31][4] ;
 wire \cur_mb_mem[31][5] ;
 wire \cur_mb_mem[31][6] ;
 wire \cur_mb_mem[31][7] ;
 wire \cur_mb_mem[32][0] ;
 wire \cur_mb_mem[32][1] ;
 wire \cur_mb_mem[32][2] ;
 wire \cur_mb_mem[32][3] ;
 wire \cur_mb_mem[32][4] ;
 wire \cur_mb_mem[32][5] ;
 wire \cur_mb_mem[32][6] ;
 wire \cur_mb_mem[32][7] ;
 wire \cur_mb_mem[33][0] ;
 wire \cur_mb_mem[33][1] ;
 wire \cur_mb_mem[33][2] ;
 wire \cur_mb_mem[33][3] ;
 wire \cur_mb_mem[33][4] ;
 wire \cur_mb_mem[33][5] ;
 wire \cur_mb_mem[33][6] ;
 wire \cur_mb_mem[33][7] ;
 wire \cur_mb_mem[34][0] ;
 wire \cur_mb_mem[34][1] ;
 wire \cur_mb_mem[34][2] ;
 wire \cur_mb_mem[34][3] ;
 wire \cur_mb_mem[34][4] ;
 wire \cur_mb_mem[34][5] ;
 wire \cur_mb_mem[34][6] ;
 wire \cur_mb_mem[34][7] ;
 wire \cur_mb_mem[35][0] ;
 wire \cur_mb_mem[35][1] ;
 wire \cur_mb_mem[35][2] ;
 wire \cur_mb_mem[35][3] ;
 wire \cur_mb_mem[35][4] ;
 wire \cur_mb_mem[35][5] ;
 wire \cur_mb_mem[35][6] ;
 wire \cur_mb_mem[35][7] ;
 wire \cur_mb_mem[36][0] ;
 wire \cur_mb_mem[36][1] ;
 wire \cur_mb_mem[36][2] ;
 wire \cur_mb_mem[36][3] ;
 wire \cur_mb_mem[36][4] ;
 wire \cur_mb_mem[36][5] ;
 wire \cur_mb_mem[36][6] ;
 wire \cur_mb_mem[36][7] ;
 wire \cur_mb_mem[37][0] ;
 wire \cur_mb_mem[37][1] ;
 wire \cur_mb_mem[37][2] ;
 wire \cur_mb_mem[37][3] ;
 wire \cur_mb_mem[37][4] ;
 wire \cur_mb_mem[37][5] ;
 wire \cur_mb_mem[37][6] ;
 wire \cur_mb_mem[37][7] ;
 wire \cur_mb_mem[38][0] ;
 wire \cur_mb_mem[38][1] ;
 wire \cur_mb_mem[38][2] ;
 wire \cur_mb_mem[38][3] ;
 wire \cur_mb_mem[38][4] ;
 wire \cur_mb_mem[38][5] ;
 wire \cur_mb_mem[38][6] ;
 wire \cur_mb_mem[38][7] ;
 wire \cur_mb_mem[39][0] ;
 wire \cur_mb_mem[39][1] ;
 wire \cur_mb_mem[39][2] ;
 wire \cur_mb_mem[39][3] ;
 wire \cur_mb_mem[39][4] ;
 wire \cur_mb_mem[39][5] ;
 wire \cur_mb_mem[39][6] ;
 wire \cur_mb_mem[39][7] ;
 wire \cur_mb_mem[3][0] ;
 wire \cur_mb_mem[3][1] ;
 wire \cur_mb_mem[3][2] ;
 wire \cur_mb_mem[3][3] ;
 wire \cur_mb_mem[3][4] ;
 wire \cur_mb_mem[3][5] ;
 wire \cur_mb_mem[3][6] ;
 wire \cur_mb_mem[3][7] ;
 wire \cur_mb_mem[40][0] ;
 wire \cur_mb_mem[40][1] ;
 wire \cur_mb_mem[40][2] ;
 wire \cur_mb_mem[40][3] ;
 wire \cur_mb_mem[40][4] ;
 wire \cur_mb_mem[40][5] ;
 wire \cur_mb_mem[40][6] ;
 wire \cur_mb_mem[40][7] ;
 wire \cur_mb_mem[41][0] ;
 wire \cur_mb_mem[41][1] ;
 wire \cur_mb_mem[41][2] ;
 wire \cur_mb_mem[41][3] ;
 wire \cur_mb_mem[41][4] ;
 wire \cur_mb_mem[41][5] ;
 wire \cur_mb_mem[41][6] ;
 wire \cur_mb_mem[41][7] ;
 wire \cur_mb_mem[42][0] ;
 wire \cur_mb_mem[42][1] ;
 wire \cur_mb_mem[42][2] ;
 wire \cur_mb_mem[42][3] ;
 wire \cur_mb_mem[42][4] ;
 wire \cur_mb_mem[42][5] ;
 wire \cur_mb_mem[42][6] ;
 wire \cur_mb_mem[42][7] ;
 wire \cur_mb_mem[43][0] ;
 wire \cur_mb_mem[43][1] ;
 wire \cur_mb_mem[43][2] ;
 wire \cur_mb_mem[43][3] ;
 wire \cur_mb_mem[43][4] ;
 wire \cur_mb_mem[43][5] ;
 wire \cur_mb_mem[43][6] ;
 wire \cur_mb_mem[43][7] ;
 wire \cur_mb_mem[44][0] ;
 wire \cur_mb_mem[44][1] ;
 wire \cur_mb_mem[44][2] ;
 wire \cur_mb_mem[44][3] ;
 wire \cur_mb_mem[44][4] ;
 wire \cur_mb_mem[44][5] ;
 wire \cur_mb_mem[44][6] ;
 wire \cur_mb_mem[44][7] ;
 wire \cur_mb_mem[45][0] ;
 wire \cur_mb_mem[45][1] ;
 wire \cur_mb_mem[45][2] ;
 wire \cur_mb_mem[45][3] ;
 wire \cur_mb_mem[45][4] ;
 wire \cur_mb_mem[45][5] ;
 wire \cur_mb_mem[45][6] ;
 wire \cur_mb_mem[45][7] ;
 wire \cur_mb_mem[46][0] ;
 wire \cur_mb_mem[46][1] ;
 wire \cur_mb_mem[46][2] ;
 wire \cur_mb_mem[46][3] ;
 wire \cur_mb_mem[46][4] ;
 wire \cur_mb_mem[46][5] ;
 wire \cur_mb_mem[46][6] ;
 wire \cur_mb_mem[46][7] ;
 wire \cur_mb_mem[47][0] ;
 wire \cur_mb_mem[47][1] ;
 wire \cur_mb_mem[47][2] ;
 wire \cur_mb_mem[47][3] ;
 wire \cur_mb_mem[47][4] ;
 wire \cur_mb_mem[47][5] ;
 wire \cur_mb_mem[47][6] ;
 wire \cur_mb_mem[47][7] ;
 wire \cur_mb_mem[48][0] ;
 wire \cur_mb_mem[48][1] ;
 wire \cur_mb_mem[48][2] ;
 wire \cur_mb_mem[48][3] ;
 wire \cur_mb_mem[48][4] ;
 wire \cur_mb_mem[48][5] ;
 wire \cur_mb_mem[48][6] ;
 wire \cur_mb_mem[48][7] ;
 wire \cur_mb_mem[49][0] ;
 wire \cur_mb_mem[49][1] ;
 wire \cur_mb_mem[49][2] ;
 wire \cur_mb_mem[49][3] ;
 wire \cur_mb_mem[49][4] ;
 wire \cur_mb_mem[49][5] ;
 wire \cur_mb_mem[49][6] ;
 wire \cur_mb_mem[49][7] ;
 wire \cur_mb_mem[4][0] ;
 wire \cur_mb_mem[4][1] ;
 wire \cur_mb_mem[4][2] ;
 wire \cur_mb_mem[4][3] ;
 wire \cur_mb_mem[4][4] ;
 wire \cur_mb_mem[4][5] ;
 wire \cur_mb_mem[4][6] ;
 wire \cur_mb_mem[4][7] ;
 wire \cur_mb_mem[50][0] ;
 wire \cur_mb_mem[50][1] ;
 wire \cur_mb_mem[50][2] ;
 wire \cur_mb_mem[50][3] ;
 wire \cur_mb_mem[50][4] ;
 wire \cur_mb_mem[50][5] ;
 wire \cur_mb_mem[50][6] ;
 wire \cur_mb_mem[50][7] ;
 wire \cur_mb_mem[51][0] ;
 wire \cur_mb_mem[51][1] ;
 wire \cur_mb_mem[51][2] ;
 wire \cur_mb_mem[51][3] ;
 wire \cur_mb_mem[51][4] ;
 wire \cur_mb_mem[51][5] ;
 wire \cur_mb_mem[51][6] ;
 wire \cur_mb_mem[51][7] ;
 wire \cur_mb_mem[52][0] ;
 wire \cur_mb_mem[52][1] ;
 wire \cur_mb_mem[52][2] ;
 wire \cur_mb_mem[52][3] ;
 wire \cur_mb_mem[52][4] ;
 wire \cur_mb_mem[52][5] ;
 wire \cur_mb_mem[52][6] ;
 wire \cur_mb_mem[52][7] ;
 wire \cur_mb_mem[53][0] ;
 wire \cur_mb_mem[53][1] ;
 wire \cur_mb_mem[53][2] ;
 wire \cur_mb_mem[53][3] ;
 wire \cur_mb_mem[53][4] ;
 wire \cur_mb_mem[53][5] ;
 wire \cur_mb_mem[53][6] ;
 wire \cur_mb_mem[53][7] ;
 wire \cur_mb_mem[54][0] ;
 wire \cur_mb_mem[54][1] ;
 wire \cur_mb_mem[54][2] ;
 wire \cur_mb_mem[54][3] ;
 wire \cur_mb_mem[54][4] ;
 wire \cur_mb_mem[54][5] ;
 wire \cur_mb_mem[54][6] ;
 wire \cur_mb_mem[54][7] ;
 wire \cur_mb_mem[55][0] ;
 wire \cur_mb_mem[55][1] ;
 wire \cur_mb_mem[55][2] ;
 wire \cur_mb_mem[55][3] ;
 wire \cur_mb_mem[55][4] ;
 wire \cur_mb_mem[55][5] ;
 wire \cur_mb_mem[55][6] ;
 wire \cur_mb_mem[55][7] ;
 wire \cur_mb_mem[56][0] ;
 wire \cur_mb_mem[56][1] ;
 wire \cur_mb_mem[56][2] ;
 wire \cur_mb_mem[56][3] ;
 wire \cur_mb_mem[56][4] ;
 wire \cur_mb_mem[56][5] ;
 wire \cur_mb_mem[56][6] ;
 wire \cur_mb_mem[56][7] ;
 wire \cur_mb_mem[57][0] ;
 wire \cur_mb_mem[57][1] ;
 wire \cur_mb_mem[57][2] ;
 wire \cur_mb_mem[57][3] ;
 wire \cur_mb_mem[57][4] ;
 wire \cur_mb_mem[57][5] ;
 wire \cur_mb_mem[57][6] ;
 wire \cur_mb_mem[57][7] ;
 wire \cur_mb_mem[58][0] ;
 wire \cur_mb_mem[58][1] ;
 wire \cur_mb_mem[58][2] ;
 wire \cur_mb_mem[58][3] ;
 wire \cur_mb_mem[58][4] ;
 wire \cur_mb_mem[58][5] ;
 wire \cur_mb_mem[58][6] ;
 wire \cur_mb_mem[58][7] ;
 wire \cur_mb_mem[59][0] ;
 wire \cur_mb_mem[59][1] ;
 wire \cur_mb_mem[59][2] ;
 wire \cur_mb_mem[59][3] ;
 wire \cur_mb_mem[59][4] ;
 wire \cur_mb_mem[59][5] ;
 wire \cur_mb_mem[59][6] ;
 wire \cur_mb_mem[59][7] ;
 wire \cur_mb_mem[5][0] ;
 wire \cur_mb_mem[5][1] ;
 wire \cur_mb_mem[5][2] ;
 wire \cur_mb_mem[5][3] ;
 wire \cur_mb_mem[5][4] ;
 wire \cur_mb_mem[5][5] ;
 wire \cur_mb_mem[5][6] ;
 wire \cur_mb_mem[5][7] ;
 wire \cur_mb_mem[60][0] ;
 wire \cur_mb_mem[60][1] ;
 wire \cur_mb_mem[60][2] ;
 wire \cur_mb_mem[60][3] ;
 wire \cur_mb_mem[60][4] ;
 wire \cur_mb_mem[60][5] ;
 wire \cur_mb_mem[60][6] ;
 wire \cur_mb_mem[60][7] ;
 wire \cur_mb_mem[61][0] ;
 wire \cur_mb_mem[61][1] ;
 wire \cur_mb_mem[61][2] ;
 wire \cur_mb_mem[61][3] ;
 wire \cur_mb_mem[61][4] ;
 wire \cur_mb_mem[61][5] ;
 wire \cur_mb_mem[61][6] ;
 wire \cur_mb_mem[61][7] ;
 wire \cur_mb_mem[62][0] ;
 wire \cur_mb_mem[62][1] ;
 wire \cur_mb_mem[62][2] ;
 wire \cur_mb_mem[62][3] ;
 wire \cur_mb_mem[62][4] ;
 wire \cur_mb_mem[62][5] ;
 wire \cur_mb_mem[62][6] ;
 wire \cur_mb_mem[62][7] ;
 wire \cur_mb_mem[63][0] ;
 wire \cur_mb_mem[63][1] ;
 wire \cur_mb_mem[63][2] ;
 wire \cur_mb_mem[63][3] ;
 wire \cur_mb_mem[63][4] ;
 wire \cur_mb_mem[63][5] ;
 wire \cur_mb_mem[63][6] ;
 wire \cur_mb_mem[63][7] ;
 wire \cur_mb_mem[64][0] ;
 wire \cur_mb_mem[64][1] ;
 wire \cur_mb_mem[64][2] ;
 wire \cur_mb_mem[64][3] ;
 wire \cur_mb_mem[64][4] ;
 wire \cur_mb_mem[64][5] ;
 wire \cur_mb_mem[64][6] ;
 wire \cur_mb_mem[64][7] ;
 wire \cur_mb_mem[65][0] ;
 wire \cur_mb_mem[65][1] ;
 wire \cur_mb_mem[65][2] ;
 wire \cur_mb_mem[65][3] ;
 wire \cur_mb_mem[65][4] ;
 wire \cur_mb_mem[65][5] ;
 wire \cur_mb_mem[65][6] ;
 wire \cur_mb_mem[65][7] ;
 wire \cur_mb_mem[66][0] ;
 wire \cur_mb_mem[66][1] ;
 wire \cur_mb_mem[66][2] ;
 wire \cur_mb_mem[66][3] ;
 wire \cur_mb_mem[66][4] ;
 wire \cur_mb_mem[66][5] ;
 wire \cur_mb_mem[66][6] ;
 wire \cur_mb_mem[66][7] ;
 wire \cur_mb_mem[67][0] ;
 wire \cur_mb_mem[67][1] ;
 wire \cur_mb_mem[67][2] ;
 wire \cur_mb_mem[67][3] ;
 wire \cur_mb_mem[67][4] ;
 wire \cur_mb_mem[67][5] ;
 wire \cur_mb_mem[67][6] ;
 wire \cur_mb_mem[67][7] ;
 wire \cur_mb_mem[68][0] ;
 wire \cur_mb_mem[68][1] ;
 wire \cur_mb_mem[68][2] ;
 wire \cur_mb_mem[68][3] ;
 wire \cur_mb_mem[68][4] ;
 wire \cur_mb_mem[68][5] ;
 wire \cur_mb_mem[68][6] ;
 wire \cur_mb_mem[68][7] ;
 wire \cur_mb_mem[69][0] ;
 wire \cur_mb_mem[69][1] ;
 wire \cur_mb_mem[69][2] ;
 wire \cur_mb_mem[69][3] ;
 wire \cur_mb_mem[69][4] ;
 wire \cur_mb_mem[69][5] ;
 wire \cur_mb_mem[69][6] ;
 wire \cur_mb_mem[69][7] ;
 wire \cur_mb_mem[6][0] ;
 wire \cur_mb_mem[6][1] ;
 wire \cur_mb_mem[6][2] ;
 wire \cur_mb_mem[6][3] ;
 wire \cur_mb_mem[6][4] ;
 wire \cur_mb_mem[6][5] ;
 wire \cur_mb_mem[6][6] ;
 wire \cur_mb_mem[6][7] ;
 wire \cur_mb_mem[70][0] ;
 wire \cur_mb_mem[70][1] ;
 wire \cur_mb_mem[70][2] ;
 wire \cur_mb_mem[70][3] ;
 wire \cur_mb_mem[70][4] ;
 wire \cur_mb_mem[70][5] ;
 wire \cur_mb_mem[70][6] ;
 wire \cur_mb_mem[70][7] ;
 wire \cur_mb_mem[71][0] ;
 wire \cur_mb_mem[71][1] ;
 wire \cur_mb_mem[71][2] ;
 wire \cur_mb_mem[71][3] ;
 wire \cur_mb_mem[71][4] ;
 wire \cur_mb_mem[71][5] ;
 wire \cur_mb_mem[71][6] ;
 wire \cur_mb_mem[71][7] ;
 wire \cur_mb_mem[72][0] ;
 wire \cur_mb_mem[72][1] ;
 wire \cur_mb_mem[72][2] ;
 wire \cur_mb_mem[72][3] ;
 wire \cur_mb_mem[72][4] ;
 wire \cur_mb_mem[72][5] ;
 wire \cur_mb_mem[72][6] ;
 wire \cur_mb_mem[72][7] ;
 wire \cur_mb_mem[73][0] ;
 wire \cur_mb_mem[73][1] ;
 wire \cur_mb_mem[73][2] ;
 wire \cur_mb_mem[73][3] ;
 wire \cur_mb_mem[73][4] ;
 wire \cur_mb_mem[73][5] ;
 wire \cur_mb_mem[73][6] ;
 wire \cur_mb_mem[73][7] ;
 wire \cur_mb_mem[74][0] ;
 wire \cur_mb_mem[74][1] ;
 wire \cur_mb_mem[74][2] ;
 wire \cur_mb_mem[74][3] ;
 wire \cur_mb_mem[74][4] ;
 wire \cur_mb_mem[74][5] ;
 wire \cur_mb_mem[74][6] ;
 wire \cur_mb_mem[74][7] ;
 wire \cur_mb_mem[75][0] ;
 wire \cur_mb_mem[75][1] ;
 wire \cur_mb_mem[75][2] ;
 wire \cur_mb_mem[75][3] ;
 wire \cur_mb_mem[75][4] ;
 wire \cur_mb_mem[75][5] ;
 wire \cur_mb_mem[75][6] ;
 wire \cur_mb_mem[75][7] ;
 wire \cur_mb_mem[76][0] ;
 wire \cur_mb_mem[76][1] ;
 wire \cur_mb_mem[76][2] ;
 wire \cur_mb_mem[76][3] ;
 wire \cur_mb_mem[76][4] ;
 wire \cur_mb_mem[76][5] ;
 wire \cur_mb_mem[76][6] ;
 wire \cur_mb_mem[76][7] ;
 wire \cur_mb_mem[77][0] ;
 wire \cur_mb_mem[77][1] ;
 wire \cur_mb_mem[77][2] ;
 wire \cur_mb_mem[77][3] ;
 wire \cur_mb_mem[77][4] ;
 wire \cur_mb_mem[77][5] ;
 wire \cur_mb_mem[77][6] ;
 wire \cur_mb_mem[77][7] ;
 wire \cur_mb_mem[78][0] ;
 wire \cur_mb_mem[78][1] ;
 wire \cur_mb_mem[78][2] ;
 wire \cur_mb_mem[78][3] ;
 wire \cur_mb_mem[78][4] ;
 wire \cur_mb_mem[78][5] ;
 wire \cur_mb_mem[78][6] ;
 wire \cur_mb_mem[78][7] ;
 wire \cur_mb_mem[79][0] ;
 wire \cur_mb_mem[79][1] ;
 wire \cur_mb_mem[79][2] ;
 wire \cur_mb_mem[79][3] ;
 wire \cur_mb_mem[79][4] ;
 wire \cur_mb_mem[79][5] ;
 wire \cur_mb_mem[79][6] ;
 wire \cur_mb_mem[79][7] ;
 wire \cur_mb_mem[7][0] ;
 wire \cur_mb_mem[7][1] ;
 wire \cur_mb_mem[7][2] ;
 wire \cur_mb_mem[7][3] ;
 wire \cur_mb_mem[7][4] ;
 wire \cur_mb_mem[7][5] ;
 wire \cur_mb_mem[7][6] ;
 wire \cur_mb_mem[7][7] ;
 wire \cur_mb_mem[80][0] ;
 wire \cur_mb_mem[80][1] ;
 wire \cur_mb_mem[80][2] ;
 wire \cur_mb_mem[80][3] ;
 wire \cur_mb_mem[80][4] ;
 wire \cur_mb_mem[80][5] ;
 wire \cur_mb_mem[80][6] ;
 wire \cur_mb_mem[80][7] ;
 wire \cur_mb_mem[81][0] ;
 wire \cur_mb_mem[81][1] ;
 wire \cur_mb_mem[81][2] ;
 wire \cur_mb_mem[81][3] ;
 wire \cur_mb_mem[81][4] ;
 wire \cur_mb_mem[81][5] ;
 wire \cur_mb_mem[81][6] ;
 wire \cur_mb_mem[81][7] ;
 wire \cur_mb_mem[82][0] ;
 wire \cur_mb_mem[82][1] ;
 wire \cur_mb_mem[82][2] ;
 wire \cur_mb_mem[82][3] ;
 wire \cur_mb_mem[82][4] ;
 wire \cur_mb_mem[82][5] ;
 wire \cur_mb_mem[82][6] ;
 wire \cur_mb_mem[82][7] ;
 wire \cur_mb_mem[83][0] ;
 wire \cur_mb_mem[83][1] ;
 wire \cur_mb_mem[83][2] ;
 wire \cur_mb_mem[83][3] ;
 wire \cur_mb_mem[83][4] ;
 wire \cur_mb_mem[83][5] ;
 wire \cur_mb_mem[83][6] ;
 wire \cur_mb_mem[83][7] ;
 wire \cur_mb_mem[84][0] ;
 wire \cur_mb_mem[84][1] ;
 wire \cur_mb_mem[84][2] ;
 wire \cur_mb_mem[84][3] ;
 wire \cur_mb_mem[84][4] ;
 wire \cur_mb_mem[84][5] ;
 wire \cur_mb_mem[84][6] ;
 wire \cur_mb_mem[84][7] ;
 wire \cur_mb_mem[85][0] ;
 wire \cur_mb_mem[85][1] ;
 wire \cur_mb_mem[85][2] ;
 wire \cur_mb_mem[85][3] ;
 wire \cur_mb_mem[85][4] ;
 wire \cur_mb_mem[85][5] ;
 wire \cur_mb_mem[85][6] ;
 wire \cur_mb_mem[85][7] ;
 wire \cur_mb_mem[86][0] ;
 wire \cur_mb_mem[86][1] ;
 wire \cur_mb_mem[86][2] ;
 wire \cur_mb_mem[86][3] ;
 wire \cur_mb_mem[86][4] ;
 wire \cur_mb_mem[86][5] ;
 wire \cur_mb_mem[86][6] ;
 wire \cur_mb_mem[86][7] ;
 wire \cur_mb_mem[87][0] ;
 wire \cur_mb_mem[87][1] ;
 wire \cur_mb_mem[87][2] ;
 wire \cur_mb_mem[87][3] ;
 wire \cur_mb_mem[87][4] ;
 wire \cur_mb_mem[87][5] ;
 wire \cur_mb_mem[87][6] ;
 wire \cur_mb_mem[87][7] ;
 wire \cur_mb_mem[88][0] ;
 wire \cur_mb_mem[88][1] ;
 wire \cur_mb_mem[88][2] ;
 wire \cur_mb_mem[88][3] ;
 wire \cur_mb_mem[88][4] ;
 wire \cur_mb_mem[88][5] ;
 wire \cur_mb_mem[88][6] ;
 wire \cur_mb_mem[88][7] ;
 wire \cur_mb_mem[89][0] ;
 wire \cur_mb_mem[89][1] ;
 wire \cur_mb_mem[89][2] ;
 wire \cur_mb_mem[89][3] ;
 wire \cur_mb_mem[89][4] ;
 wire \cur_mb_mem[89][5] ;
 wire \cur_mb_mem[89][6] ;
 wire \cur_mb_mem[89][7] ;
 wire \cur_mb_mem[8][0] ;
 wire \cur_mb_mem[8][1] ;
 wire \cur_mb_mem[8][2] ;
 wire \cur_mb_mem[8][3] ;
 wire \cur_mb_mem[8][4] ;
 wire \cur_mb_mem[8][5] ;
 wire \cur_mb_mem[8][6] ;
 wire \cur_mb_mem[8][7] ;
 wire \cur_mb_mem[90][0] ;
 wire \cur_mb_mem[90][1] ;
 wire \cur_mb_mem[90][2] ;
 wire \cur_mb_mem[90][3] ;
 wire \cur_mb_mem[90][4] ;
 wire \cur_mb_mem[90][5] ;
 wire \cur_mb_mem[90][6] ;
 wire \cur_mb_mem[90][7] ;
 wire \cur_mb_mem[91][0] ;
 wire \cur_mb_mem[91][1] ;
 wire \cur_mb_mem[91][2] ;
 wire \cur_mb_mem[91][3] ;
 wire \cur_mb_mem[91][4] ;
 wire \cur_mb_mem[91][5] ;
 wire \cur_mb_mem[91][6] ;
 wire \cur_mb_mem[91][7] ;
 wire \cur_mb_mem[92][0] ;
 wire \cur_mb_mem[92][1] ;
 wire \cur_mb_mem[92][2] ;
 wire \cur_mb_mem[92][3] ;
 wire \cur_mb_mem[92][4] ;
 wire \cur_mb_mem[92][5] ;
 wire \cur_mb_mem[92][6] ;
 wire \cur_mb_mem[92][7] ;
 wire \cur_mb_mem[93][0] ;
 wire \cur_mb_mem[93][1] ;
 wire \cur_mb_mem[93][2] ;
 wire \cur_mb_mem[93][3] ;
 wire \cur_mb_mem[93][4] ;
 wire \cur_mb_mem[93][5] ;
 wire \cur_mb_mem[93][6] ;
 wire \cur_mb_mem[93][7] ;
 wire \cur_mb_mem[94][0] ;
 wire \cur_mb_mem[94][1] ;
 wire \cur_mb_mem[94][2] ;
 wire \cur_mb_mem[94][3] ;
 wire \cur_mb_mem[94][4] ;
 wire \cur_mb_mem[94][5] ;
 wire \cur_mb_mem[94][6] ;
 wire \cur_mb_mem[94][7] ;
 wire \cur_mb_mem[95][0] ;
 wire \cur_mb_mem[95][1] ;
 wire \cur_mb_mem[95][2] ;
 wire \cur_mb_mem[95][3] ;
 wire \cur_mb_mem[95][4] ;
 wire \cur_mb_mem[95][5] ;
 wire \cur_mb_mem[95][6] ;
 wire \cur_mb_mem[95][7] ;
 wire \cur_mb_mem[96][0] ;
 wire \cur_mb_mem[96][1] ;
 wire \cur_mb_mem[96][2] ;
 wire \cur_mb_mem[96][3] ;
 wire \cur_mb_mem[96][4] ;
 wire \cur_mb_mem[96][5] ;
 wire \cur_mb_mem[96][6] ;
 wire \cur_mb_mem[96][7] ;
 wire \cur_mb_mem[97][0] ;
 wire \cur_mb_mem[97][1] ;
 wire \cur_mb_mem[97][2] ;
 wire \cur_mb_mem[97][3] ;
 wire \cur_mb_mem[97][4] ;
 wire \cur_mb_mem[97][5] ;
 wire \cur_mb_mem[97][6] ;
 wire \cur_mb_mem[97][7] ;
 wire \cur_mb_mem[98][0] ;
 wire \cur_mb_mem[98][1] ;
 wire \cur_mb_mem[98][2] ;
 wire \cur_mb_mem[98][3] ;
 wire \cur_mb_mem[98][4] ;
 wire \cur_mb_mem[98][5] ;
 wire \cur_mb_mem[98][6] ;
 wire \cur_mb_mem[98][7] ;
 wire \cur_mb_mem[99][0] ;
 wire \cur_mb_mem[99][1] ;
 wire \cur_mb_mem[99][2] ;
 wire \cur_mb_mem[99][3] ;
 wire \cur_mb_mem[99][4] ;
 wire \cur_mb_mem[99][5] ;
 wire \cur_mb_mem[99][6] ;
 wire \cur_mb_mem[99][7] ;
 wire \cur_mb_mem[9][0] ;
 wire \cur_mb_mem[9][1] ;
 wire \cur_mb_mem[9][2] ;
 wire \cur_mb_mem[9][3] ;
 wire \cur_mb_mem[9][4] ;
 wire \cur_mb_mem[9][5] ;
 wire \cur_mb_mem[9][6] ;
 wire \cur_mb_mem[9][7] ;
 wire \current_accum_sad[0] ;
 wire \current_accum_sad[10] ;
 wire \current_accum_sad[11] ;
 wire \current_accum_sad[12] ;
 wire \current_accum_sad[13] ;
 wire \current_accum_sad[14] ;
 wire \current_accum_sad[15] ;
 wire \current_accum_sad[1] ;
 wire \current_accum_sad[2] ;
 wire \current_accum_sad[3] ;
 wire \current_accum_sad[4] ;
 wire \current_accum_sad[5] ;
 wire \current_accum_sad[6] ;
 wire \current_accum_sad[7] ;
 wire \current_accum_sad[8] ;
 wire \current_accum_sad[9] ;
 wire \min_sad_reg[0] ;
 wire \min_sad_reg[10] ;
 wire \min_sad_reg[11] ;
 wire \min_sad_reg[12] ;
 wire \min_sad_reg[13] ;
 wire \min_sad_reg[14] ;
 wire \min_sad_reg[15] ;
 wire \min_sad_reg[1] ;
 wire \min_sad_reg[2] ;
 wire \min_sad_reg[3] ;
 wire \min_sad_reg[4] ;
 wire \min_sad_reg[5] ;
 wire \min_sad_reg[6] ;
 wire \min_sad_reg[7] ;
 wire \min_sad_reg[8] ;
 wire \min_sad_reg[9] ;
 wire \pixel_cnt[0] ;
 wire \pixel_cnt[1] ;
 wire \pixel_cnt[2] ;
 wire \pixel_cnt[3] ;
 wire \pixel_cnt[4] ;
 wire \pixel_cnt[5] ;
 wire \pixel_cnt[6] ;
 wire \pixel_cnt[7] ;
 wire \pixel_cnt[8] ;
 wire \point_cnt[0] ;
 wire \point_cnt[1] ;
 wire \point_cnt[2] ;
 wire \point_cnt[3] ;
 wire \shex_center_x[0] ;
 wire \shex_center_x[1] ;
 wire \shex_center_x[2] ;
 wire \shex_center_x[3] ;
 wire \shex_center_x[4] ;
 wire \shex_center_x[5] ;
 wire \shex_center_x[6] ;
 wire \shex_center_y[0] ;
 wire \shex_center_y[1] ;
 wire \shex_center_y[2] ;
 wire \shex_center_y[3] ;
 wire \shex_center_y[4] ;
 wire \shex_center_y[5] ;
 wire \shex_center_y[6] ;
 wire shex_load;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[6] ;
 wire \state[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_316_clk;
 wire clknet_leaf_317_clk;
 wire clknet_leaf_318_clk;
 wire clknet_leaf_319_clk;
 wire clknet_leaf_320_clk;
 wire clknet_leaf_321_clk;
 wire clknet_leaf_322_clk;
 wire clknet_leaf_323_clk;
 wire clknet_leaf_324_clk;
 wire clknet_leaf_325_clk;
 wire clknet_leaf_326_clk;
 wire clknet_leaf_327_clk;
 wire clknet_leaf_328_clk;
 wire clknet_leaf_329_clk;
 wire clknet_leaf_330_clk;
 wire clknet_leaf_331_clk;
 wire clknet_leaf_332_clk;
 wire clknet_leaf_333_clk;
 wire clknet_leaf_334_clk;
 wire clknet_leaf_335_clk;
 wire clknet_leaf_336_clk;
 wire clknet_leaf_337_clk;
 wire clknet_leaf_338_clk;
 wire clknet_leaf_339_clk;
 wire clknet_leaf_340_clk;
 wire clknet_leaf_341_clk;
 wire clknet_leaf_342_clk;
 wire clknet_leaf_343_clk;
 wire clknet_leaf_344_clk;
 wire clknet_leaf_345_clk;
 wire clknet_leaf_346_clk;
 wire clknet_leaf_347_clk;
 wire clknet_leaf_348_clk;
 wire clknet_leaf_349_clk;
 wire clknet_leaf_350_clk;
 wire clknet_leaf_351_clk;
 wire clknet_leaf_352_clk;
 wire clknet_leaf_353_clk;
 wire clknet_leaf_354_clk;
 wire clknet_leaf_355_clk;
 wire clknet_leaf_356_clk;
 wire clknet_leaf_357_clk;
 wire clknet_leaf_358_clk;
 wire clknet_leaf_359_clk;
 wire clknet_leaf_360_clk;
 wire clknet_leaf_361_clk;
 wire clknet_leaf_362_clk;
 wire clknet_leaf_363_clk;
 wire clknet_leaf_364_clk;
 wire clknet_leaf_365_clk;
 wire clknet_leaf_366_clk;
 wire clknet_leaf_367_clk;
 wire clknet_leaf_368_clk;
 wire clknet_leaf_369_clk;
 wire clknet_leaf_370_clk;
 wire clknet_leaf_371_clk;
 wire clknet_leaf_372_clk;
 wire clknet_leaf_373_clk;
 wire clknet_leaf_374_clk;
 wire clknet_leaf_375_clk;
 wire clknet_leaf_376_clk;
 wire clknet_leaf_377_clk;
 wire clknet_leaf_378_clk;
 wire clknet_leaf_379_clk;
 wire clknet_leaf_380_clk;
 wire clknet_leaf_381_clk;
 wire clknet_leaf_382_clk;
 wire clknet_leaf_383_clk;
 wire clknet_leaf_384_clk;
 wire clknet_leaf_385_clk;
 wire clknet_leaf_386_clk;
 wire clknet_leaf_387_clk;
 wire clknet_leaf_388_clk;
 wire clknet_leaf_389_clk;
 wire clknet_leaf_390_clk;
 wire clknet_leaf_391_clk;
 wire clknet_leaf_392_clk;
 wire clknet_leaf_393_clk;
 wire clknet_leaf_394_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;

 sky130_fd_sc_hd__buf_2 _09335_ (.A(\pixel_cnt[1] ),
    .X(_04420_));
 sky130_fd_sc_hd__buf_2 _09336_ (.A(\pixel_cnt[0] ),
    .X(_04421_));
 sky130_fd_sc_hd__and4_2 _09337_ (.A(_04420_),
    .B(_04421_),
    .C(\pixel_cnt[2] ),
    .D(\pixel_cnt[3] ),
    .X(_04422_));
 sky130_fd_sc_hd__buf_4 _09338_ (.A(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__buf_8 _09339_ (.A(_04423_),
    .X(_04424_));
 sky130_fd_sc_hd__clkbuf_4 _09340_ (.A(\pixel_cnt[4] ),
    .X(_04425_));
 sky130_fd_sc_hd__clkbuf_4 _09341_ (.A(\pixel_cnt[5] ),
    .X(_04426_));
 sky130_fd_sc_hd__clkbuf_4 _09342_ (.A(\pixel_cnt[7] ),
    .X(_04427_));
 sky130_fd_sc_hd__clkbuf_4 _09343_ (.A(\pixel_cnt[6] ),
    .X(_04428_));
 sky130_fd_sc_hd__and4_4 _09344_ (.A(_04425_),
    .B(_04426_),
    .C(_04427_),
    .D(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__buf_8 _09345_ (.A(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__clkbuf_8 _09346_ (.A(_04430_),
    .X(_04431_));
 sky130_fd_sc_hd__clkbuf_16 _09347_ (.A(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__nand2_4 _09348_ (.A(_04424_),
    .B(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__nor2_1 _09349_ (.A(\pixel_cnt[8] ),
    .B(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__buf_2 _09350_ (.A(\point_cnt[2] ),
    .X(_04435_));
 sky130_fd_sc_hd__buf_2 _09351_ (.A(\point_cnt[0] ),
    .X(_04436_));
 sky130_fd_sc_hd__clkbuf_4 _09352_ (.A(\point_cnt[1] ),
    .X(_04437_));
 sky130_fd_sc_hd__and2b_1 _09353_ (.A_N(_04436_),
    .B(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__clkbuf_4 _09354_ (.A(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__and3b_1 _09355_ (.A_N(\point_cnt[3] ),
    .B(_04435_),
    .C(_04439_),
    .X(_04440_));
 sky130_fd_sc_hd__and3_1 _09356_ (.A(\state[6] ),
    .B(_04434_),
    .C(_04440_),
    .X(_04441_));
 sky130_fd_sc_hd__buf_1 _09357_ (.A(_04441_),
    .X(_00001_));
 sky130_fd_sc_hd__or2_2 _09358_ (.A(\pixel_cnt[8] ),
    .B(_04433_),
    .X(_04442_));
 sky130_fd_sc_hd__clkbuf_8 _09359_ (.A(\state[4] ),
    .X(_04443_));
 sky130_fd_sc_hd__buf_8 _09360_ (.A(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__a22o_1 _09361_ (.A1(net1786),
    .A2(net138),
    .B1(_04442_),
    .B2(_04444_),
    .X(_00005_));
 sky130_fd_sc_hd__inv_2 _09362_ (.A(\state[1] ),
    .Y(_04445_));
 sky130_fd_sc_hd__or4_1 _09363_ (.A(\best_point_idx[1] ),
    .B(\best_point_idx[0] ),
    .C(\best_point_idx[3] ),
    .D(net291),
    .X(_04446_));
 sky130_fd_sc_hd__nor2_1 _09364_ (.A(_04445_),
    .B(net292),
    .Y(_00002_));
 sky130_fd_sc_hd__clkbuf_4 _09365_ (.A(\state[6] ),
    .X(_04447_));
 sky130_fd_sc_hd__nand2_1 _09366_ (.A(_04434_),
    .B(_04440_),
    .Y(_04448_));
 sky130_fd_sc_hd__a21o_1 _09367_ (.A1(_04447_),
    .A2(_04448_),
    .B1(net389),
    .X(_00006_));
 sky130_fd_sc_hd__buf_4 _09368_ (.A(\state[7] ),
    .X(_04449_));
 sky130_fd_sc_hd__nand2_2 _09369_ (.A(_04437_),
    .B(\point_cnt[0] ),
    .Y(_04450_));
 sky130_fd_sc_hd__nor3_1 _09370_ (.A(\point_cnt[3] ),
    .B(_04435_),
    .C(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__or3b_1 _09371_ (.A(shex_load),
    .B(_04442_),
    .C_N(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__inv_2 _09372_ (.A(\state[3] ),
    .Y(_04453_));
 sky130_fd_sc_hd__o2bb2ai_1 _09373_ (.A1_N(_04449_),
    .A2_N(net138),
    .B1(_04452_),
    .B2(_04453_),
    .Y(_00007_));
 sky130_fd_sc_hd__clkbuf_4 _09374_ (.A(\state[3] ),
    .X(_04454_));
 sky130_fd_sc_hd__a21o_1 _09375_ (.A1(_04454_),
    .A2(_04452_),
    .B1(net310),
    .X(_00004_));
 sky130_fd_sc_hd__clkbuf_4 _09376_ (.A(\state[1] ),
    .X(_04455_));
 sky130_fd_sc_hd__a22o_1 _09377_ (.A1(_04444_),
    .A2(_04434_),
    .B1(net292),
    .B2(_04455_),
    .X(_00003_));
 sky130_fd_sc_hd__nand2_1 _09378_ (.A(net33),
    .B(net1),
    .Y(_04456_));
 sky130_fd_sc_hd__or2_1 _09379_ (.A(net33),
    .B(net1),
    .X(_04457_));
 sky130_fd_sc_hd__buf_2 _09380_ (.A(\pixel_cnt[0] ),
    .X(_04458_));
 sky130_fd_sc_hd__buf_4 _09381_ (.A(_04458_),
    .X(_04459_));
 sky130_fd_sc_hd__a21o_1 _09382_ (.A1(_04456_),
    .A2(_04457_),
    .B1(_04459_),
    .X(_04460_));
 sky130_fd_sc_hd__nand3_1 _09383_ (.A(_04459_),
    .B(_04456_),
    .C(_04457_),
    .Y(_04461_));
 sky130_fd_sc_hd__or2_1 _09384_ (.A(\state[6] ),
    .B(\state[3] ),
    .X(_04462_));
 sky130_fd_sc_hd__clkbuf_8 _09385_ (.A(_04462_),
    .X(_04463_));
 sky130_fd_sc_hd__clkbuf_8 _09386_ (.A(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__and2_1 _09387_ (.A(_04459_),
    .B(net105),
    .X(_04465_));
 sky130_fd_sc_hd__nor2_1 _09388_ (.A(_04459_),
    .B(net105),
    .Y(_04466_));
 sky130_fd_sc_hd__nor2_1 _09389_ (.A(_04465_),
    .B(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__nand2_1 _09390_ (.A(\cand_x[0] ),
    .B(net33),
    .Y(_04468_));
 sky130_fd_sc_hd__or2_1 _09391_ (.A(\cand_x[0] ),
    .B(net33),
    .X(_04469_));
 sky130_fd_sc_hd__and2_1 _09392_ (.A(_04468_),
    .B(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__buf_4 _09393_ (.A(\cand_x[6] ),
    .X(_04471_));
 sky130_fd_sc_hd__clkbuf_4 _09394_ (.A(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__buf_4 _09395_ (.A(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__clkbuf_4 _09396_ (.A(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__buf_6 _09397_ (.A(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__or2_1 _09398_ (.A(_04475_),
    .B(net56),
    .X(_04476_));
 sky130_fd_sc_hd__nand2_1 _09399_ (.A(_04475_),
    .B(net56),
    .Y(_04477_));
 sky130_fd_sc_hd__nand2_2 _09400_ (.A(_04476_),
    .B(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__or2_2 _09401_ (.A(\cand_x[5] ),
    .B(net60),
    .X(_04479_));
 sky130_fd_sc_hd__or2_1 _09402_ (.A(\cand_x[4] ),
    .B(net59),
    .X(_04480_));
 sky130_fd_sc_hd__nor2_1 _09403_ (.A(\cand_x[3] ),
    .B(net58),
    .Y(_04481_));
 sky130_fd_sc_hd__nor2_1 _09404_ (.A(\cand_x[2] ),
    .B(net55),
    .Y(_04482_));
 sky130_fd_sc_hd__nor2_1 _09405_ (.A(\cand_x[1] ),
    .B(net44),
    .Y(_04483_));
 sky130_fd_sc_hd__nand2_1 _09406_ (.A(\cand_x[1] ),
    .B(net44),
    .Y(_04484_));
 sky130_fd_sc_hd__o21a_1 _09407_ (.A1(_04468_),
    .A2(_04483_),
    .B1(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__nand2_1 _09408_ (.A(\cand_x[2] ),
    .B(net55),
    .Y(_04486_));
 sky130_fd_sc_hd__o21a_1 _09409_ (.A1(_04482_),
    .A2(_04485_),
    .B1(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__and2_1 _09410_ (.A(\cand_x[3] ),
    .B(net58),
    .X(_04488_));
 sky130_fd_sc_hd__o21bai_2 _09411_ (.A1(_04481_),
    .A2(_04487_),
    .B1_N(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__and2_1 _09412_ (.A(\cand_x[4] ),
    .B(net59),
    .X(_04490_));
 sky130_fd_sc_hd__a221o_2 _09413_ (.A1(\cand_x[5] ),
    .A2(net60),
    .B1(_04480_),
    .B2(_04489_),
    .C1(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__xor2_2 _09414_ (.A(_04471_),
    .B(net62),
    .X(_04492_));
 sky130_fd_sc_hd__xor2_2 _09415_ (.A(_04471_),
    .B(net61),
    .X(_04493_));
 sky130_fd_sc_hd__and2_1 _09416_ (.A(_04492_),
    .B(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__buf_4 _09417_ (.A(_04471_),
    .X(_04495_));
 sky130_fd_sc_hd__o21a_1 _09418_ (.A1(net62),
    .A2(net61),
    .B1(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__a31o_2 _09419_ (.A1(_04479_),
    .A2(_04491_),
    .A3(_04494_),
    .B1(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__xor2_1 _09420_ (.A(_04472_),
    .B(net35),
    .X(_04498_));
 sky130_fd_sc_hd__and2_1 _09421_ (.A(_04471_),
    .B(net34),
    .X(_04499_));
 sky130_fd_sc_hd__nor2_1 _09422_ (.A(_04472_),
    .B(net34),
    .Y(_04500_));
 sky130_fd_sc_hd__nor2_1 _09423_ (.A(_04499_),
    .B(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__xor2_2 _09424_ (.A(_04472_),
    .B(net64),
    .X(_04502_));
 sky130_fd_sc_hd__and2_1 _09425_ (.A(_04471_),
    .B(net63),
    .X(_04503_));
 sky130_fd_sc_hd__nor2_1 _09426_ (.A(_04472_),
    .B(net63),
    .Y(_04504_));
 sky130_fd_sc_hd__nor2_2 _09427_ (.A(_04503_),
    .B(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__and4_1 _09428_ (.A(_04498_),
    .B(_04501_),
    .C(_04502_),
    .D(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__xor2_1 _09429_ (.A(_04495_),
    .B(net37),
    .X(_04507_));
 sky130_fd_sc_hd__and2_1 _09430_ (.A(_04471_),
    .B(net36),
    .X(_04508_));
 sky130_fd_sc_hd__nor2_1 _09431_ (.A(_04472_),
    .B(net36),
    .Y(_04509_));
 sky130_fd_sc_hd__nor2_1 _09432_ (.A(_04508_),
    .B(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__and2_1 _09433_ (.A(_04471_),
    .B(net38),
    .X(_04511_));
 sky130_fd_sc_hd__nor2_1 _09434_ (.A(_04472_),
    .B(net38),
    .Y(_04512_));
 sky130_fd_sc_hd__nor2_1 _09435_ (.A(_04511_),
    .B(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__xor2_1 _09436_ (.A(_04495_),
    .B(net39),
    .X(_04514_));
 sky130_fd_sc_hd__and4_1 _09437_ (.A(_04507_),
    .B(_04510_),
    .C(_04513_),
    .D(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__nand3_2 _09438_ (.A(_04497_),
    .B(_04506_),
    .C(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__o21a_1 _09439_ (.A1(net64),
    .A2(net63),
    .B1(_04472_),
    .X(_04517_));
 sky130_fd_sc_hd__a211o_1 _09440_ (.A1(_04473_),
    .A2(net35),
    .B1(_04499_),
    .C1(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__o21a_1 _09441_ (.A1(net37),
    .A2(net36),
    .B1(_04473_),
    .X(_04519_));
 sky130_fd_sc_hd__a2111oi_4 _09442_ (.A1(_04473_),
    .A2(net39),
    .B1(_04511_),
    .C1(_04518_),
    .D1(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__xnor2_1 _09443_ (.A(_04495_),
    .B(net43),
    .Y(_04521_));
 sky130_fd_sc_hd__nand2_1 _09444_ (.A(_04495_),
    .B(net42),
    .Y(_04522_));
 sky130_fd_sc_hd__or2_1 _09445_ (.A(_04472_),
    .B(net42),
    .X(_04523_));
 sky130_fd_sc_hd__nand2_1 _09446_ (.A(_04522_),
    .B(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__xnor2_2 _09447_ (.A(_04495_),
    .B(net41),
    .Y(_04525_));
 sky130_fd_sc_hd__nand2_1 _09448_ (.A(_04495_),
    .B(net40),
    .Y(_04526_));
 sky130_fd_sc_hd__or2_1 _09449_ (.A(_04472_),
    .B(net40),
    .X(_04527_));
 sky130_fd_sc_hd__nand2_1 _09450_ (.A(_04526_),
    .B(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__or4_1 _09451_ (.A(_04521_),
    .B(_04524_),
    .C(_04525_),
    .D(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__xnor2_2 _09452_ (.A(_04495_),
    .B(net46),
    .Y(_04530_));
 sky130_fd_sc_hd__nand2_1 _09453_ (.A(_04471_),
    .B(net45),
    .Y(_04531_));
 sky130_fd_sc_hd__or2_1 _09454_ (.A(_04471_),
    .B(net45),
    .X(_04532_));
 sky130_fd_sc_hd__and2_1 _09455_ (.A(_04531_),
    .B(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__inv_2 _09456_ (.A(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2_1 _09457_ (.A(_04495_),
    .B(net47),
    .Y(_04535_));
 sky130_fd_sc_hd__or2_1 _09458_ (.A(_04495_),
    .B(net47),
    .X(_04536_));
 sky130_fd_sc_hd__nand2_1 _09459_ (.A(_04535_),
    .B(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__xnor2_1 _09460_ (.A(_04473_),
    .B(net48),
    .Y(_04538_));
 sky130_fd_sc_hd__or4_1 _09461_ (.A(_04530_),
    .B(_04534_),
    .C(_04537_),
    .D(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__a211o_1 _09462_ (.A1(_04516_),
    .A2(_04520_),
    .B1(_04529_),
    .C1(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__o41a_1 _09463_ (.A1(net43),
    .A2(net42),
    .A3(net41),
    .A4(net40),
    .B1(_04474_),
    .X(_04541_));
 sky130_fd_sc_hd__o41a_1 _09464_ (.A1(net48),
    .A2(net47),
    .A3(net46),
    .A4(net45),
    .B1(_04474_),
    .X(_04542_));
 sky130_fd_sc_hd__nor2_1 _09465_ (.A(_04541_),
    .B(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__xnor2_1 _09466_ (.A(_04473_),
    .B(net50),
    .Y(_04544_));
 sky130_fd_sc_hd__nand2_1 _09467_ (.A(_04474_),
    .B(net49),
    .Y(_04545_));
 sky130_fd_sc_hd__or2_1 _09468_ (.A(_04473_),
    .B(net49),
    .X(_04546_));
 sky130_fd_sc_hd__nand2_1 _09469_ (.A(_04545_),
    .B(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__or2_1 _09470_ (.A(_04544_),
    .B(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__xnor2_1 _09471_ (.A(_04474_),
    .B(net52),
    .Y(_04549_));
 sky130_fd_sc_hd__nand2_1 _09472_ (.A(_04473_),
    .B(net51),
    .Y(_04550_));
 sky130_fd_sc_hd__or2_1 _09473_ (.A(_04473_),
    .B(net51),
    .X(_04551_));
 sky130_fd_sc_hd__and2_1 _09474_ (.A(_04550_),
    .B(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__inv_2 _09475_ (.A(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__a2111oi_1 _09476_ (.A1(_04540_),
    .A2(_04543_),
    .B1(_04548_),
    .C1(_04549_),
    .D1(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__o41a_1 _09477_ (.A1(net52),
    .A2(net51),
    .A3(net50),
    .A4(net49),
    .B1(_04475_),
    .X(_04555_));
 sky130_fd_sc_hd__nand2_1 _09478_ (.A(_04474_),
    .B(net53),
    .Y(_04556_));
 sky130_fd_sc_hd__or2_1 _09479_ (.A(_04474_),
    .B(net53),
    .X(_04557_));
 sky130_fd_sc_hd__and2_1 _09480_ (.A(_04556_),
    .B(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__o21ai_1 _09481_ (.A1(net212),
    .A2(_04555_),
    .B1(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__nor2_1 _09482_ (.A(_04475_),
    .B(net54),
    .Y(_04560_));
 sky130_fd_sc_hd__nand2_1 _09483_ (.A(_04475_),
    .B(net54),
    .Y(_04561_));
 sky130_fd_sc_hd__o211a_1 _09484_ (.A1(_04559_),
    .A2(_04560_),
    .B1(_04561_),
    .C1(_04556_),
    .X(_04562_));
 sky130_fd_sc_hd__xnor2_1 _09485_ (.A(_04478_),
    .B(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__or2b_1 _09486_ (.A(_04560_),
    .B_N(_04561_),
    .X(_04564_));
 sky130_fd_sc_hd__nand2_1 _09487_ (.A(_04556_),
    .B(_04559_),
    .Y(_04565_));
 sky130_fd_sc_hd__xor2_1 _09488_ (.A(_04564_),
    .B(_04565_),
    .X(_04566_));
 sky130_fd_sc_hd__o21a_1 _09489_ (.A1(net46),
    .A2(net45),
    .B1(_04474_),
    .X(_04567_));
 sky130_fd_sc_hd__a21oi_1 _09490_ (.A1(_04516_),
    .A2(_04520_),
    .B1(_04529_),
    .Y(_04568_));
 sky130_fd_sc_hd__inv_2 _09491_ (.A(_04530_),
    .Y(_04569_));
 sky130_fd_sc_hd__o211a_1 _09492_ (.A1(_04568_),
    .A2(_04541_),
    .B1(_04533_),
    .C1(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__o21bai_1 _09493_ (.A1(_04567_),
    .A2(_04570_),
    .B1_N(_04537_),
    .Y(_04571_));
 sky130_fd_sc_hd__a21oi_1 _09494_ (.A1(_04535_),
    .A2(_04571_),
    .B1(_04538_),
    .Y(_04572_));
 sky130_fd_sc_hd__and3_1 _09495_ (.A(_04535_),
    .B(_04538_),
    .C(_04571_),
    .X(_04573_));
 sky130_fd_sc_hd__or3b_1 _09496_ (.A(_04567_),
    .B(_04570_),
    .C_N(_04537_),
    .X(_04574_));
 sky130_fd_sc_hd__nand2_1 _09497_ (.A(_04516_),
    .B(_04520_),
    .Y(_04575_));
 sky130_fd_sc_hd__a21bo_1 _09498_ (.A1(_04575_),
    .A2(_04527_),
    .B1_N(_04526_),
    .X(_04576_));
 sky130_fd_sc_hd__xnor2_1 _09499_ (.A(_04525_),
    .B(_04576_),
    .Y(_04577_));
 sky130_fd_sc_hd__a21oi_1 _09500_ (.A1(_04497_),
    .A2(_04505_),
    .B1(_04503_),
    .Y(_04578_));
 sky130_fd_sc_hd__xnor2_1 _09501_ (.A(_04502_),
    .B(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__xnor2_2 _09502_ (.A(_04497_),
    .B(_04505_),
    .Y(_04580_));
 sky130_fd_sc_hd__nand2_1 _09503_ (.A(_04479_),
    .B(_04491_),
    .Y(_04581_));
 sky130_fd_sc_hd__xor2_2 _09504_ (.A(_04581_),
    .B(_04493_),
    .X(_04582_));
 sky130_fd_sc_hd__and2b_1 _09505_ (.A_N(_04490_),
    .B(_04480_),
    .X(_04583_));
 sky130_fd_sc_hd__xnor2_1 _09506_ (.A(_04583_),
    .B(_04489_),
    .Y(_04584_));
 sky130_fd_sc_hd__inv_2 _09507_ (.A(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__nor2_1 _09508_ (.A(_04488_),
    .B(_04481_),
    .Y(_04586_));
 sky130_fd_sc_hd__xnor2_1 _09509_ (.A(_04487_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__or2_1 _09510_ (.A(\cand_x[1] ),
    .B(net44),
    .X(_04588_));
 sky130_fd_sc_hd__nand2_1 _09511_ (.A(_04484_),
    .B(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__xor2_2 _09512_ (.A(_04468_),
    .B(_04589_),
    .X(_04590_));
 sky130_fd_sc_hd__and2b_1 _09513_ (.A_N(_04482_),
    .B(_04486_),
    .X(_04591_));
 sky130_fd_sc_hd__xnor2_1 _09514_ (.A(_04485_),
    .B(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__or4_1 _09515_ (.A(_04470_),
    .B(_04587_),
    .C(_04590_),
    .D(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__nand2_1 _09516_ (.A(\cand_x[5] ),
    .B(net60),
    .Y(_04594_));
 sky130_fd_sc_hd__nand2_1 _09517_ (.A(_04479_),
    .B(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__a21o_1 _09518_ (.A1(_04480_),
    .A2(_04489_),
    .B1(_04490_),
    .X(_04596_));
 sky130_fd_sc_hd__xnor2_2 _09519_ (.A(_04595_),
    .B(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__a21oi_2 _09520_ (.A1(_04585_),
    .A2(_04593_),
    .B1(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__a32o_1 _09521_ (.A1(_04479_),
    .A2(_04491_),
    .A3(_04493_),
    .B1(net61),
    .B2(_04473_),
    .X(_04599_));
 sky130_fd_sc_hd__xor2_2 _09522_ (.A(_04492_),
    .B(_04599_),
    .X(_04600_));
 sky130_fd_sc_hd__o21ba_1 _09523_ (.A1(_04582_),
    .A2(_04598_),
    .B1_N(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__a21o_1 _09524_ (.A1(_04497_),
    .A2(_04506_),
    .B1(_04518_),
    .X(_04602_));
 sky130_fd_sc_hd__xnor2_1 _09525_ (.A(_04510_),
    .B(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__o21ai_1 _09526_ (.A1(_04580_),
    .A2(_04601_),
    .B1(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__xnor2_1 _09527_ (.A(_04575_),
    .B(_04528_),
    .Y(_04605_));
 sky130_fd_sc_hd__a31o_1 _09528_ (.A1(_04497_),
    .A2(_04502_),
    .A3(_04505_),
    .B1(_04517_),
    .X(_04606_));
 sky130_fd_sc_hd__xor2_1 _09529_ (.A(_04501_),
    .B(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__or4_1 _09530_ (.A(_04579_),
    .B(_04604_),
    .C(_04605_),
    .D(_04607_),
    .X(_04608_));
 sky130_fd_sc_hd__o21ai_1 _09531_ (.A1(_04568_),
    .A2(_04541_),
    .B1(_04533_),
    .Y(_04609_));
 sky130_fd_sc_hd__or3_1 _09532_ (.A(_04568_),
    .B(_04533_),
    .C(_04541_),
    .X(_04610_));
 sky130_fd_sc_hd__o21ai_1 _09533_ (.A1(net41),
    .A2(net40),
    .B1(_04474_),
    .Y(_04611_));
 sky130_fd_sc_hd__a211o_1 _09534_ (.A1(_04516_),
    .A2(_04520_),
    .B1(_04525_),
    .C1(_04528_),
    .X(_04612_));
 sky130_fd_sc_hd__nand3_1 _09535_ (.A(_04524_),
    .B(_04611_),
    .C(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__a21o_1 _09536_ (.A1(_04611_),
    .A2(_04612_),
    .B1(_04524_),
    .X(_04614_));
 sky130_fd_sc_hd__a22o_1 _09537_ (.A1(_04609_),
    .A2(_04610_),
    .B1(_04613_),
    .B2(_04614_),
    .X(_04615_));
 sky130_fd_sc_hd__a2111oi_1 _09538_ (.A1(_04571_),
    .A2(_04574_),
    .B1(_04577_),
    .C1(_04608_),
    .D1(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__a21oi_1 _09539_ (.A1(_04522_),
    .A2(_04614_),
    .B1(_04521_),
    .Y(_04617_));
 sky130_fd_sc_hd__and3_1 _09540_ (.A(_04521_),
    .B(_04522_),
    .C(_04614_),
    .X(_04618_));
 sky130_fd_sc_hd__a21oi_1 _09541_ (.A1(_04531_),
    .A2(_04609_),
    .B1(_04530_),
    .Y(_04619_));
 sky130_fd_sc_hd__and3_1 _09542_ (.A(_04530_),
    .B(_04531_),
    .C(_04609_),
    .X(_04620_));
 sky130_fd_sc_hd__o22a_1 _09543_ (.A1(_04617_),
    .A2(_04618_),
    .B1(_04619_),
    .B2(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__o211a_1 _09544_ (.A1(_04572_),
    .A2(_04573_),
    .B1(_04616_),
    .C1(_04621_),
    .X(_04622_));
 sky130_fd_sc_hd__a21oi_1 _09545_ (.A1(_04540_),
    .A2(_04543_),
    .B1(_04548_),
    .Y(_04623_));
 sky130_fd_sc_hd__o21a_1 _09546_ (.A1(net50),
    .A2(net49),
    .B1(_04474_),
    .X(_04624_));
 sky130_fd_sc_hd__o21ai_1 _09547_ (.A1(_04623_),
    .A2(_04624_),
    .B1(_04552_),
    .Y(_04625_));
 sky130_fd_sc_hd__a21oi_1 _09548_ (.A1(_04550_),
    .A2(_04625_),
    .B1(_04549_),
    .Y(_04626_));
 sky130_fd_sc_hd__and3_1 _09549_ (.A(_04549_),
    .B(_04550_),
    .C(_04625_),
    .X(_04627_));
 sky130_fd_sc_hd__nand2_1 _09550_ (.A(_04540_),
    .B(_04543_),
    .Y(_04628_));
 sky130_fd_sc_hd__a21bo_1 _09551_ (.A1(_04628_),
    .A2(_04546_),
    .B1_N(_04545_),
    .X(_04629_));
 sky130_fd_sc_hd__xor2_1 _09552_ (.A(_04544_),
    .B(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__or3_1 _09553_ (.A(_04558_),
    .B(net213),
    .C(_04555_),
    .X(_04631_));
 sky130_fd_sc_hd__nand2_1 _09554_ (.A(_04559_),
    .B(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__or3_1 _09555_ (.A(_04623_),
    .B(_04552_),
    .C(_04624_),
    .X(_04633_));
 sky130_fd_sc_hd__xnor2_1 _09556_ (.A(_04628_),
    .B(_04547_),
    .Y(_04634_));
 sky130_fd_sc_hd__a21oi_1 _09557_ (.A1(_04501_),
    .A2(_04606_),
    .B1(_04499_),
    .Y(_04635_));
 sky130_fd_sc_hd__xnor2_1 _09558_ (.A(_04498_),
    .B(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__a31o_1 _09559_ (.A1(_04507_),
    .A2(_04510_),
    .A3(_04602_),
    .B1(_04519_),
    .X(_04637_));
 sky130_fd_sc_hd__xor2_1 _09560_ (.A(_04513_),
    .B(_04637_),
    .X(_04638_));
 sky130_fd_sc_hd__a21oi_1 _09561_ (.A1(_04510_),
    .A2(_04602_),
    .B1(_04508_),
    .Y(_04639_));
 sky130_fd_sc_hd__xnor2_1 _09562_ (.A(_04507_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__or3_1 _09563_ (.A(_04636_),
    .B(_04638_),
    .C(_04640_),
    .X(_04641_));
 sky130_fd_sc_hd__a21oi_1 _09564_ (.A1(_04513_),
    .A2(_04637_),
    .B1(_04511_),
    .Y(_04642_));
 sky130_fd_sc_hd__xnor2_1 _09565_ (.A(_04514_),
    .B(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hd__a2111oi_1 _09566_ (.A1(_04625_),
    .A2(_04633_),
    .B1(_04634_),
    .C1(_04641_),
    .D1(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__o2111a_1 _09567_ (.A1(_04626_),
    .A2(_04627_),
    .B1(_04630_),
    .C1(_04632_),
    .D1(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__and4_4 _09568_ (.A(_04563_),
    .B(_04566_),
    .C(_04622_),
    .D(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__o21ai_4 _09569_ (.A1(_04478_),
    .A2(_04562_),
    .B1(_04477_),
    .Y(_04647_));
 sky130_fd_sc_hd__xor2_4 _09570_ (.A(_04475_),
    .B(net57),
    .X(_04648_));
 sky130_fd_sc_hd__xnor2_4 _09571_ (.A(_04647_),
    .B(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__and2_1 _09572_ (.A(_04646_),
    .B(_04649_),
    .X(_04650_));
 sky130_fd_sc_hd__nand2_1 _09573_ (.A(_04470_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__xnor2_1 _09574_ (.A(_04467_),
    .B(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__a32o_2 _09575_ (.A1(_04444_),
    .A2(_04460_),
    .A3(_04461_),
    .B1(_04464_),
    .B2(_04652_),
    .X(net140));
 sky130_fd_sc_hd__buf_2 _09576_ (.A(\pixel_cnt[1] ),
    .X(_04653_));
 sky130_fd_sc_hd__buf_4 _09577_ (.A(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__nor2_1 _09578_ (.A(_04654_),
    .B(net116),
    .Y(_04655_));
 sky130_fd_sc_hd__and2_1 _09579_ (.A(_04654_),
    .B(net116),
    .X(_04656_));
 sky130_fd_sc_hd__nor2_1 _09580_ (.A(_04655_),
    .B(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__nand2_1 _09581_ (.A(_04590_),
    .B(_04650_),
    .Y(_04658_));
 sky130_fd_sc_hd__xnor2_2 _09582_ (.A(_04657_),
    .B(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__a31o_1 _09583_ (.A1(_04467_),
    .A2(_04470_),
    .A3(_04650_),
    .B1(_04465_),
    .X(_04660_));
 sky130_fd_sc_hd__nor2_1 _09584_ (.A(_04659_),
    .B(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__nand2_1 _09585_ (.A(_04659_),
    .B(_04660_),
    .Y(_04662_));
 sky130_fd_sc_hd__nand2_1 _09586_ (.A(_04463_),
    .B(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__xor2_2 _09587_ (.A(net44),
    .B(net12),
    .X(_04664_));
 sky130_fd_sc_hd__xnor2_1 _09588_ (.A(_04654_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__a21o_1 _09589_ (.A1(_04456_),
    .A2(_04461_),
    .B1(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__nand2_1 _09590_ (.A(_04443_),
    .B(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__a31o_1 _09591_ (.A1(_04456_),
    .A2(_04461_),
    .A3(_04665_),
    .B1(_04667_),
    .X(_04668_));
 sky130_fd_sc_hd__o21ai_4 _09592_ (.A1(_04661_),
    .A2(_04663_),
    .B1(_04668_),
    .Y(net151));
 sky130_fd_sc_hd__buf_2 _09593_ (.A(\pixel_cnt[2] ),
    .X(_04669_));
 sky130_fd_sc_hd__buf_4 _09594_ (.A(_04669_),
    .X(_04670_));
 sky130_fd_sc_hd__xor2_1 _09595_ (.A(net55),
    .B(net23),
    .X(_04671_));
 sky130_fd_sc_hd__xnor2_1 _09596_ (.A(_04670_),
    .B(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__and2_1 _09597_ (.A(net44),
    .B(net12),
    .X(_04673_));
 sky130_fd_sc_hd__a21oi_2 _09598_ (.A1(_04654_),
    .A2(_04664_),
    .B1(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__xnor2_1 _09599_ (.A(_04672_),
    .B(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__nand2_1 _09600_ (.A(_04666_),
    .B(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__or2_1 _09601_ (.A(_04666_),
    .B(_04675_),
    .X(_04677_));
 sky130_fd_sc_hd__nor2_1 _09602_ (.A(_04670_),
    .B(net127),
    .Y(_04678_));
 sky130_fd_sc_hd__and2_1 _09603_ (.A(_04670_),
    .B(net127),
    .X(_04679_));
 sky130_fd_sc_hd__nor2_1 _09604_ (.A(_04678_),
    .B(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__and3_1 _09605_ (.A(_04592_),
    .B(_04646_),
    .C(_04649_),
    .X(_04681_));
 sky130_fd_sc_hd__xnor2_1 _09606_ (.A(_04680_),
    .B(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__a31o_1 _09607_ (.A1(_04590_),
    .A2(_04650_),
    .A3(_04657_),
    .B1(_04656_),
    .X(_04683_));
 sky130_fd_sc_hd__xnor2_1 _09608_ (.A(_04682_),
    .B(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__xnor2_1 _09609_ (.A(_04662_),
    .B(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__a32o_2 _09610_ (.A1(_04444_),
    .A2(_04676_),
    .A3(_04677_),
    .B1(_04685_),
    .B2(_04464_),
    .X(net162));
 sky130_fd_sc_hd__nor2_4 _09611_ (.A(\state[6] ),
    .B(\state[3] ),
    .Y(_04686_));
 sky130_fd_sc_hd__clkbuf_8 _09612_ (.A(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__buf_6 _09613_ (.A(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__buf_4 _09614_ (.A(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__and2b_1 _09615_ (.A_N(_04682_),
    .B(_04683_),
    .X(_04690_));
 sky130_fd_sc_hd__buf_2 _09616_ (.A(\pixel_cnt[3] ),
    .X(_04691_));
 sky130_fd_sc_hd__clkbuf_4 _09617_ (.A(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__or2_1 _09618_ (.A(_04692_),
    .B(net130),
    .X(_04693_));
 sky130_fd_sc_hd__nand2_1 _09619_ (.A(_04692_),
    .B(net130),
    .Y(_04694_));
 sky130_fd_sc_hd__nand2_1 _09620_ (.A(_04693_),
    .B(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__and3_1 _09621_ (.A(_04587_),
    .B(_04646_),
    .C(_04649_),
    .X(_04696_));
 sky130_fd_sc_hd__xor2_2 _09622_ (.A(_04695_),
    .B(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__a21o_1 _09623_ (.A1(_04680_),
    .A2(_04681_),
    .B1(_04679_),
    .X(_04698_));
 sky130_fd_sc_hd__xnor2_2 _09624_ (.A(_04697_),
    .B(_04698_),
    .Y(_04699_));
 sky130_fd_sc_hd__and2_1 _09625_ (.A(_04690_),
    .B(_04699_),
    .X(_04700_));
 sky130_fd_sc_hd__nor2_1 _09626_ (.A(_04690_),
    .B(_04699_),
    .Y(_04701_));
 sky130_fd_sc_hd__or2_1 _09627_ (.A(_04700_),
    .B(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__and3_1 _09628_ (.A(_04659_),
    .B(_04660_),
    .C(_04684_),
    .X(_04703_));
 sky130_fd_sc_hd__mux2_1 _09629_ (.A0(_04702_),
    .A1(_04699_),
    .S(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__xor2_1 _09630_ (.A(net58),
    .B(net26),
    .X(_04705_));
 sky130_fd_sc_hd__xnor2_1 _09631_ (.A(_04692_),
    .B(_04705_),
    .Y(_04706_));
 sky130_fd_sc_hd__and2_1 _09632_ (.A(net55),
    .B(net23),
    .X(_04707_));
 sky130_fd_sc_hd__a21oi_1 _09633_ (.A1(_04670_),
    .A2(_04671_),
    .B1(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__xnor2_1 _09634_ (.A(_04706_),
    .B(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__or3_1 _09635_ (.A(_04672_),
    .B(_04674_),
    .C(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__o21ai_1 _09636_ (.A1(_04672_),
    .A2(_04674_),
    .B1(_04709_),
    .Y(_04711_));
 sky130_fd_sc_hd__nand2_1 _09637_ (.A(_04710_),
    .B(_04711_),
    .Y(_04712_));
 sky130_fd_sc_hd__or3_1 _09638_ (.A(_04666_),
    .B(_04675_),
    .C(_04709_),
    .X(_04713_));
 sky130_fd_sc_hd__a21boi_1 _09639_ (.A1(_04677_),
    .A2(_04712_),
    .B1_N(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__a2bb2o_4 _09640_ (.A1_N(_04689_),
    .A2_N(_04704_),
    .B1(_04714_),
    .B2(_04444_),
    .X(net165));
 sky130_fd_sc_hd__nor2_1 _09641_ (.A(_04706_),
    .B(_04708_),
    .Y(_04715_));
 sky130_fd_sc_hd__nand2_1 _09642_ (.A(net59),
    .B(net27),
    .Y(_04716_));
 sky130_fd_sc_hd__or2_1 _09643_ (.A(net59),
    .B(net27),
    .X(_04717_));
 sky130_fd_sc_hd__nand2_1 _09644_ (.A(_04716_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__and2_1 _09645_ (.A(net58),
    .B(net26),
    .X(_04719_));
 sky130_fd_sc_hd__a21o_1 _09646_ (.A1(_04692_),
    .A2(_04705_),
    .B1(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__xnor2_1 _09647_ (.A(_04718_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__xnor2_1 _09648_ (.A(_04715_),
    .B(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__and3_1 _09649_ (.A(_04710_),
    .B(_04713_),
    .C(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__buf_4 _09650_ (.A(_04443_),
    .X(_04724_));
 sky130_fd_sc_hd__a21o_1 _09651_ (.A1(_04710_),
    .A2(_04713_),
    .B1(_04722_),
    .X(_04725_));
 sky130_fd_sc_hd__nand2_1 _09652_ (.A(_04724_),
    .B(_04725_),
    .Y(_04726_));
 sky130_fd_sc_hd__and4_1 _09653_ (.A(_04659_),
    .B(_04660_),
    .C(_04684_),
    .D(_04699_),
    .X(_04727_));
 sky130_fd_sc_hd__or2b_1 _09654_ (.A(_04697_),
    .B_N(_04698_),
    .X(_04728_));
 sky130_fd_sc_hd__inv_2 _09655_ (.A(net131),
    .Y(_04729_));
 sky130_fd_sc_hd__a21bo_1 _09656_ (.A1(_04584_),
    .A2(_04646_),
    .B1_N(_04649_),
    .X(_04730_));
 sky130_fd_sc_hd__xnor2_1 _09657_ (.A(_04729_),
    .B(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__a21bo_1 _09658_ (.A1(_04693_),
    .A2(_04696_),
    .B1_N(_04694_),
    .X(_04732_));
 sky130_fd_sc_hd__xor2_1 _09659_ (.A(_04731_),
    .B(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__xor2_1 _09660_ (.A(_04728_),
    .B(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__o21ai_2 _09661_ (.A1(_04700_),
    .A2(_04727_),
    .B1(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__o31a_1 _09662_ (.A1(_04700_),
    .A2(_04727_),
    .A3(_04734_),
    .B1(_04463_),
    .X(_04736_));
 sky130_fd_sc_hd__a2bb2o_4 _09663_ (.A1_N(_04723_),
    .A2_N(_04726_),
    .B1(_04735_),
    .B2(_04736_),
    .X(net166));
 sky130_fd_sc_hd__and2b_1 _09664_ (.A_N(_04731_),
    .B(_04732_),
    .X(_04737_));
 sky130_fd_sc_hd__clkbuf_4 _09665_ (.A(_04425_),
    .X(_04738_));
 sky130_fd_sc_hd__inv_2 _09666_ (.A(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__nor2_1 _09667_ (.A(_04729_),
    .B(_04730_),
    .Y(_04740_));
 sky130_fd_sc_hd__buf_6 _09668_ (.A(net65),
    .X(_04741_));
 sky130_fd_sc_hd__nand2_2 _09669_ (.A(\cand_y[0] ),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__or2_1 _09670_ (.A(\cand_y[0] ),
    .B(_04741_),
    .X(_04743_));
 sky130_fd_sc_hd__nand2_4 _09671_ (.A(_04742_),
    .B(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__clkbuf_4 _09672_ (.A(\cand_y[6] ),
    .X(_04745_));
 sky130_fd_sc_hd__clkbuf_4 _09673_ (.A(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__clkbuf_4 _09674_ (.A(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__clkbuf_4 _09675_ (.A(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__nand2_1 _09676_ (.A(_04748_),
    .B(net81),
    .Y(_04749_));
 sky130_fd_sc_hd__or2_1 _09677_ (.A(_04748_),
    .B(net81),
    .X(_04750_));
 sky130_fd_sc_hd__nand2_1 _09678_ (.A(_04749_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__inv_2 _09679_ (.A(_04745_),
    .Y(_04752_));
 sky130_fd_sc_hd__inv_2 _09680_ (.A(net77),
    .Y(_04753_));
 sky130_fd_sc_hd__nor2_1 _09681_ (.A(_04752_),
    .B(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__nor2_1 _09682_ (.A(_04746_),
    .B(net77),
    .Y(_04755_));
 sky130_fd_sc_hd__nor2_1 _09683_ (.A(_04754_),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__xor2_1 _09684_ (.A(_04747_),
    .B(net78),
    .X(_04757_));
 sky130_fd_sc_hd__and2_1 _09685_ (.A(_04756_),
    .B(_04757_),
    .X(_04758_));
 sky130_fd_sc_hd__inv_2 _09686_ (.A(net79),
    .Y(_04759_));
 sky130_fd_sc_hd__nor2_1 _09687_ (.A(_04752_),
    .B(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__buf_4 _09688_ (.A(_04747_),
    .X(_04761_));
 sky130_fd_sc_hd__nor2_1 _09689_ (.A(_04761_),
    .B(net79),
    .Y(_04762_));
 sky130_fd_sc_hd__nor2_1 _09690_ (.A(_04760_),
    .B(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__xor2_2 _09691_ (.A(_04761_),
    .B(net80),
    .X(_04764_));
 sky130_fd_sc_hd__and3_1 _09692_ (.A(_04758_),
    .B(_04763_),
    .C(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__inv_2 _09693_ (.A(net72),
    .Y(_04766_));
 sky130_fd_sc_hd__nor2_1 _09694_ (.A(_04752_),
    .B(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hd__nor2_1 _09695_ (.A(_04746_),
    .B(net72),
    .Y(_04768_));
 sky130_fd_sc_hd__nor2_1 _09696_ (.A(_04767_),
    .B(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__buf_4 _09697_ (.A(net73),
    .X(_04770_));
 sky130_fd_sc_hd__xor2_1 _09698_ (.A(_04746_),
    .B(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__and2_1 _09699_ (.A(_04769_),
    .B(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__clkbuf_4 _09700_ (.A(net75),
    .X(_04773_));
 sky130_fd_sc_hd__xor2_1 _09701_ (.A(_04747_),
    .B(_04773_),
    .X(_04774_));
 sky130_fd_sc_hd__inv_2 _09702_ (.A(net74),
    .Y(_04775_));
 sky130_fd_sc_hd__nor2_1 _09703_ (.A(_04752_),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__nor2_1 _09704_ (.A(_04747_),
    .B(net74),
    .Y(_04777_));
 sky130_fd_sc_hd__nor2_1 _09705_ (.A(_04776_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__and3_1 _09706_ (.A(_04772_),
    .B(_04774_),
    .C(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__buf_6 _09707_ (.A(net94),
    .X(_04780_));
 sky130_fd_sc_hd__buf_6 _09708_ (.A(net93),
    .X(_04781_));
 sky130_fd_sc_hd__o21ai_1 _09709_ (.A1(_04780_),
    .A2(_04781_),
    .B1(_04747_),
    .Y(_04782_));
 sky130_fd_sc_hd__nor2_1 _09710_ (.A(\cand_y[3] ),
    .B(net90),
    .Y(_04783_));
 sky130_fd_sc_hd__buf_6 _09711_ (.A(net87),
    .X(_04784_));
 sky130_fd_sc_hd__nand2_2 _09712_ (.A(\cand_y[2] ),
    .B(_04784_),
    .Y(_04785_));
 sky130_fd_sc_hd__or2_1 _09713_ (.A(\cand_y[2] ),
    .B(net87),
    .X(_04786_));
 sky130_fd_sc_hd__nand2_4 _09714_ (.A(_04785_),
    .B(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__buf_6 _09715_ (.A(net76),
    .X(_04788_));
 sky130_fd_sc_hd__nor2_1 _09716_ (.A(\cand_y[1] ),
    .B(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__nand2_1 _09717_ (.A(\cand_y[1] ),
    .B(_04788_),
    .Y(_04790_));
 sky130_fd_sc_hd__o21a_2 _09718_ (.A1(_04742_),
    .A2(_04789_),
    .B1(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__nand2_1 _09719_ (.A(\cand_y[3] ),
    .B(net90),
    .Y(_04792_));
 sky130_fd_sc_hd__o211a_1 _09720_ (.A1(_04787_),
    .A2(_04791_),
    .B1(_04792_),
    .C1(_04785_),
    .X(_04793_));
 sky130_fd_sc_hd__xor2_1 _09721_ (.A(_04745_),
    .B(_04781_),
    .X(_04794_));
 sky130_fd_sc_hd__xor2_1 _09722_ (.A(_04745_),
    .B(_04780_),
    .X(_04795_));
 sky130_fd_sc_hd__nand2_1 _09723_ (.A(_04794_),
    .B(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__nand2_1 _09724_ (.A(\cand_y[4] ),
    .B(net91),
    .Y(_04797_));
 sky130_fd_sc_hd__or2_1 _09725_ (.A(\cand_y[4] ),
    .B(net91),
    .X(_04798_));
 sky130_fd_sc_hd__nand2_1 _09726_ (.A(_04797_),
    .B(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__nand2_1 _09727_ (.A(\cand_y[5] ),
    .B(net92),
    .Y(_04800_));
 sky130_fd_sc_hd__or2_1 _09728_ (.A(\cand_y[5] ),
    .B(net92),
    .X(_04801_));
 sky130_fd_sc_hd__nand2_2 _09729_ (.A(_04800_),
    .B(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__or3_1 _09730_ (.A(_04796_),
    .B(_04799_),
    .C(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__a21bo_1 _09731_ (.A1(_04797_),
    .A2(_04800_),
    .B1_N(_04801_),
    .X(_04804_));
 sky130_fd_sc_hd__or2_1 _09732_ (.A(_04796_),
    .B(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__o31a_1 _09733_ (.A1(_04783_),
    .A2(_04793_),
    .A3(_04803_),
    .B1(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__buf_4 _09734_ (.A(net95),
    .X(_04807_));
 sky130_fd_sc_hd__xor2_1 _09735_ (.A(_04745_),
    .B(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__or2_1 _09736_ (.A(_04745_),
    .B(net96),
    .X(_04809_));
 sky130_fd_sc_hd__clkbuf_4 _09737_ (.A(net96),
    .X(_04810_));
 sky130_fd_sc_hd__nand2_1 _09738_ (.A(_04745_),
    .B(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__and3_1 _09739_ (.A(_04808_),
    .B(_04809_),
    .C(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__inv_2 _09740_ (.A(_04812_),
    .Y(_04813_));
 sky130_fd_sc_hd__clkbuf_4 _09741_ (.A(net67),
    .X(_04814_));
 sky130_fd_sc_hd__xnor2_1 _09742_ (.A(_04746_),
    .B(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand2_1 _09743_ (.A(_04746_),
    .B(net66),
    .Y(_04816_));
 sky130_fd_sc_hd__or2_1 _09744_ (.A(_04745_),
    .B(net66),
    .X(_04817_));
 sky130_fd_sc_hd__nand2_1 _09745_ (.A(_04816_),
    .B(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__a2111oi_1 _09746_ (.A1(_04782_),
    .A2(_04806_),
    .B1(_04813_),
    .C1(_04815_),
    .D1(_04818_),
    .Y(_04819_));
 sky130_fd_sc_hd__or2_1 _09747_ (.A(_04745_),
    .B(net69),
    .X(_04820_));
 sky130_fd_sc_hd__nand2_1 _09748_ (.A(_04746_),
    .B(net69),
    .Y(_04821_));
 sky130_fd_sc_hd__nand2_1 _09749_ (.A(_04820_),
    .B(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__nand2_1 _09750_ (.A(_04746_),
    .B(net68),
    .Y(_04823_));
 sky130_fd_sc_hd__or2_1 _09751_ (.A(_04745_),
    .B(net68),
    .X(_04824_));
 sky130_fd_sc_hd__and2_1 _09752_ (.A(_04823_),
    .B(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__buf_4 _09753_ (.A(net71),
    .X(_04826_));
 sky130_fd_sc_hd__xor2_1 _09754_ (.A(_04746_),
    .B(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__inv_2 _09755_ (.A(net70),
    .Y(_04828_));
 sky130_fd_sc_hd__nor2_1 _09756_ (.A(_04752_),
    .B(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__nor2_1 _09757_ (.A(_04746_),
    .B(net70),
    .Y(_04830_));
 sky130_fd_sc_hd__nor2_1 _09758_ (.A(_04829_),
    .B(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__and4b_1 _09759_ (.A_N(_04822_),
    .B(_04825_),
    .C(_04827_),
    .D(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__o41a_1 _09760_ (.A1(_04814_),
    .A2(net66),
    .A3(_04810_),
    .A4(_04807_),
    .B1(_04747_),
    .X(_04833_));
 sky130_fd_sc_hd__o41a_1 _09761_ (.A1(_04826_),
    .A2(net70),
    .A3(net69),
    .A4(net68),
    .B1(_04761_),
    .X(_04834_));
 sky130_fd_sc_hd__a211o_2 _09762_ (.A1(net219),
    .A2(_04832_),
    .B1(_04833_),
    .C1(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__o41a_1 _09763_ (.A1(_04773_),
    .A2(net74),
    .A3(_04770_),
    .A4(net72),
    .B1(_04761_),
    .X(_04836_));
 sky130_fd_sc_hd__o41a_1 _09764_ (.A1(net80),
    .A2(net79),
    .A3(net78),
    .A4(net77),
    .B1(_04761_),
    .X(_04837_));
 sky130_fd_sc_hd__or2_1 _09765_ (.A(_04836_),
    .B(_04837_),
    .X(_04838_));
 sky130_fd_sc_hd__a31o_1 _09766_ (.A1(_04765_),
    .A2(_04779_),
    .A3(net288),
    .B1(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__or2b_1 _09767_ (.A(_04751_),
    .B_N(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__xor2_1 _09768_ (.A(_04748_),
    .B(net82),
    .X(_04841_));
 sky130_fd_sc_hd__a21oi_1 _09769_ (.A1(_04749_),
    .A2(_04840_),
    .B1(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__o21ai_1 _09770_ (.A1(net219),
    .A2(_04833_),
    .B1(_04825_),
    .Y(_04843_));
 sky130_fd_sc_hd__nand2_1 _09771_ (.A(_04823_),
    .B(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hd__xnor2_1 _09772_ (.A(_04822_),
    .B(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__nand2_1 _09773_ (.A(_04782_),
    .B(_04806_),
    .Y(_04846_));
 sky130_fd_sc_hd__o21a_1 _09774_ (.A1(_04810_),
    .A2(_04807_),
    .B1(_04761_),
    .X(_04847_));
 sky130_fd_sc_hd__a21oi_1 _09775_ (.A1(_04846_),
    .A2(_04812_),
    .B1(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__o21ai_1 _09776_ (.A1(_04818_),
    .A2(_04848_),
    .B1(_04816_),
    .Y(_04849_));
 sky130_fd_sc_hd__xnor2_1 _09777_ (.A(_04815_),
    .B(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__clkbuf_8 _09778_ (.A(_04748_),
    .X(_04851_));
 sky130_fd_sc_hd__a21o_1 _09779_ (.A1(_04779_),
    .A2(net289),
    .B1(_04836_),
    .X(_04852_));
 sky130_fd_sc_hd__a221o_1 _09780_ (.A1(_04851_),
    .A2(net78),
    .B1(_04758_),
    .B2(_04852_),
    .C1(_04754_),
    .X(_04853_));
 sky130_fd_sc_hd__a21oi_1 _09781_ (.A1(_04763_),
    .A2(_04853_),
    .B1(_04760_),
    .Y(_04854_));
 sky130_fd_sc_hd__a32o_1 _09782_ (.A1(_04841_),
    .A2(_04749_),
    .A3(_04840_),
    .B1(_04854_),
    .B2(_04764_),
    .X(_04855_));
 sky130_fd_sc_hd__or4_4 _09783_ (.A(_04842_),
    .B(_04845_),
    .C(_04850_),
    .D(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__or2_1 _09784_ (.A(_04851_),
    .B(net88),
    .X(_04857_));
 sky130_fd_sc_hd__nand2_1 _09785_ (.A(_04851_),
    .B(net88),
    .Y(_04858_));
 sky130_fd_sc_hd__nand2_1 _09786_ (.A(_04857_),
    .B(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__and2_1 _09787_ (.A(_04748_),
    .B(net85),
    .X(_04860_));
 sky130_fd_sc_hd__nor2_1 _09788_ (.A(_04761_),
    .B(net85),
    .Y(_04861_));
 sky130_fd_sc_hd__nor2_1 _09789_ (.A(_04860_),
    .B(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__and3_1 _09790_ (.A(_04841_),
    .B(_04749_),
    .C(_04750_),
    .X(_04863_));
 sky130_fd_sc_hd__nand2_1 _09791_ (.A(_04761_),
    .B(net84),
    .Y(_04864_));
 sky130_fd_sc_hd__or2_1 _09792_ (.A(_04747_),
    .B(net84),
    .X(_04865_));
 sky130_fd_sc_hd__o211a_1 _09793_ (.A1(_04748_),
    .A2(net83),
    .B1(_04864_),
    .C1(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__o41a_1 _09794_ (.A1(net84),
    .A2(net83),
    .A3(net82),
    .A4(net81),
    .B1(_04748_),
    .X(_04867_));
 sky130_fd_sc_hd__a31o_1 _09795_ (.A1(_04839_),
    .A2(_04863_),
    .A3(_04866_),
    .B1(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__or2_1 _09796_ (.A(_04747_),
    .B(net86),
    .X(_04869_));
 sky130_fd_sc_hd__o21a_1 _09797_ (.A1(net86),
    .A2(net85),
    .B1(_04851_),
    .X(_04870_));
 sky130_fd_sc_hd__a31o_1 _09798_ (.A1(_04862_),
    .A2(_04868_),
    .A3(_04869_),
    .B1(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__xnor2_1 _09799_ (.A(_04859_),
    .B(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__nor2_1 _09800_ (.A(_04764_),
    .B(_04854_),
    .Y(_04873_));
 sky130_fd_sc_hd__xor2_1 _09801_ (.A(_04851_),
    .B(net83),
    .X(_04874_));
 sky130_fd_sc_hd__o21a_1 _09802_ (.A1(net82),
    .A2(net81),
    .B1(_04851_),
    .X(_04875_));
 sky130_fd_sc_hd__a21oi_1 _09803_ (.A1(_04839_),
    .A2(_04863_),
    .B1(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__xnor2_1 _09804_ (.A(_04874_),
    .B(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__xor2_1 _09805_ (.A(_04862_),
    .B(_04868_),
    .X(_04878_));
 sky130_fd_sc_hd__xor2_1 _09806_ (.A(_04763_),
    .B(_04853_),
    .X(_04879_));
 sky130_fd_sc_hd__o211a_1 _09807_ (.A1(_04822_),
    .A2(_04843_),
    .B1(_04823_),
    .C1(_04821_),
    .X(_04880_));
 sky130_fd_sc_hd__o21ba_1 _09808_ (.A1(_04830_),
    .A2(_04880_),
    .B1_N(_04829_),
    .X(_04881_));
 sky130_fd_sc_hd__xnor2_1 _09809_ (.A(_04827_),
    .B(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__or4_1 _09810_ (.A(_04877_),
    .B(_04878_),
    .C(_04879_),
    .D(_04882_),
    .X(_04883_));
 sky130_fd_sc_hd__a221o_1 _09811_ (.A1(_04748_),
    .A2(_04770_),
    .B1(_04772_),
    .B2(_04835_),
    .C1(_04767_),
    .X(_04884_));
 sky130_fd_sc_hd__nand2_1 _09812_ (.A(_04778_),
    .B(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__or2_1 _09813_ (.A(_04778_),
    .B(_04884_),
    .X(_04886_));
 sky130_fd_sc_hd__xor2_1 _09814_ (.A(_04756_),
    .B(_04852_),
    .X(_04887_));
 sky130_fd_sc_hd__xnor2_1 _09815_ (.A(_04839_),
    .B(_04751_),
    .Y(_04888_));
 sky130_fd_sc_hd__a211o_1 _09816_ (.A1(_04885_),
    .A2(_04886_),
    .B1(_04887_),
    .C1(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__xnor2_1 _09817_ (.A(_04831_),
    .B(_04880_),
    .Y(_04890_));
 sky130_fd_sc_hd__a21oi_1 _09818_ (.A1(_04769_),
    .A2(_04835_),
    .B1(_04767_),
    .Y(_04891_));
 sky130_fd_sc_hd__xnor2_1 _09819_ (.A(_04771_),
    .B(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__or3_1 _09820_ (.A(net286),
    .B(_04825_),
    .C(_04833_),
    .X(_04893_));
 sky130_fd_sc_hd__xor2_1 _09821_ (.A(_04818_),
    .B(_04848_),
    .X(_04894_));
 sky130_fd_sc_hd__nor2_1 _09822_ (.A(_04747_),
    .B(_04781_),
    .Y(_04895_));
 sky130_fd_sc_hd__o41a_1 _09823_ (.A1(_04783_),
    .A2(_04793_),
    .A3(_04799_),
    .A4(_04802_),
    .B1(_04804_),
    .X(_04896_));
 sky130_fd_sc_hd__nand2_1 _09824_ (.A(_04761_),
    .B(_04781_),
    .Y(_04897_));
 sky130_fd_sc_hd__o21ai_1 _09825_ (.A1(_04895_),
    .A2(_04896_),
    .B1(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__xnor2_2 _09826_ (.A(net282),
    .B(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__xnor2_1 _09827_ (.A(net290),
    .B(_04896_),
    .Y(_04900_));
 sky130_fd_sc_hd__inv_2 _09828_ (.A(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__o31a_1 _09829_ (.A1(_04783_),
    .A2(_04793_),
    .A3(_04799_),
    .B1(_04797_),
    .X(_04902_));
 sky130_fd_sc_hd__xor2_2 _09830_ (.A(_04802_),
    .B(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__inv_2 _09831_ (.A(_04903_),
    .Y(_04904_));
 sky130_fd_sc_hd__or2_1 _09832_ (.A(_04783_),
    .B(_04793_),
    .X(_04905_));
 sky130_fd_sc_hd__xnor2_1 _09833_ (.A(_04905_),
    .B(_04799_),
    .Y(_04906_));
 sky130_fd_sc_hd__xor2_1 _09834_ (.A(_04787_),
    .B(_04791_),
    .X(_04907_));
 sky130_fd_sc_hd__or2_1 _09835_ (.A(\cand_y[1] ),
    .B(_04788_),
    .X(_04908_));
 sky130_fd_sc_hd__nand2_1 _09836_ (.A(_04790_),
    .B(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__xnor2_2 _09837_ (.A(_04742_),
    .B(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__inv_2 _09838_ (.A(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__nor2_1 _09839_ (.A(_04907_),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__o21ai_1 _09840_ (.A1(_04787_),
    .A2(_04791_),
    .B1(_04785_),
    .Y(_04913_));
 sky130_fd_sc_hd__and2b_1 _09841_ (.A_N(_04783_),
    .B(_04792_),
    .X(_04914_));
 sky130_fd_sc_hd__xnor2_1 _09842_ (.A(_04913_),
    .B(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__and4_1 _09843_ (.A(_04744_),
    .B(_04906_),
    .C(_04912_),
    .D(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__nor4_1 _09844_ (.A(_04899_),
    .B(_04901_),
    .C(_04904_),
    .D(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__a211o_1 _09845_ (.A1(_04843_),
    .A2(_04893_),
    .B1(_04894_),
    .C1(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__xor2_1 _09846_ (.A(_04769_),
    .B(_04835_),
    .X(_04919_));
 sky130_fd_sc_hd__nand2_1 _09847_ (.A(_04846_),
    .B(_04812_),
    .Y(_04920_));
 sky130_fd_sc_hd__o31a_1 _09848_ (.A1(_04810_),
    .A2(_04846_),
    .A3(_04808_),
    .B1(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__nor3_1 _09849_ (.A(_04748_),
    .B(net84),
    .C(net83),
    .Y(_04922_));
 sky130_fd_sc_hd__nor3_1 _09850_ (.A(_04748_),
    .B(net86),
    .C(net85),
    .Y(_04923_));
 sky130_fd_sc_hd__nand2_1 _09851_ (.A(_04761_),
    .B(net86),
    .Y(_04924_));
 sky130_fd_sc_hd__and3b_1 _09852_ (.A_N(_04861_),
    .B(_04869_),
    .C(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__o22a_1 _09853_ (.A1(_04866_),
    .A2(_04922_),
    .B1(_04923_),
    .B2(_04925_),
    .X(_04926_));
 sky130_fd_sc_hd__or3b_1 _09854_ (.A(_04919_),
    .B(_04921_),
    .C_N(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__or4_1 _09855_ (.A(_04890_),
    .B(_04892_),
    .C(_04918_),
    .D(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__a21oi_1 _09856_ (.A1(_04778_),
    .A2(_04884_),
    .B1(_04776_),
    .Y(_04929_));
 sky130_fd_sc_hd__xnor2_1 _09857_ (.A(_04774_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__a21oi_1 _09858_ (.A1(_04756_),
    .A2(_04852_),
    .B1(_04754_),
    .Y(_04931_));
 sky130_fd_sc_hd__xnor2_1 _09859_ (.A(_04757_),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__or4_1 _09860_ (.A(_04889_),
    .B(_04928_),
    .C(_04930_),
    .D(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__or4_4 _09861_ (.A(_04872_),
    .B(_04873_),
    .C(_04883_),
    .D(_04933_),
    .X(_04934_));
 sky130_fd_sc_hd__a21bo_2 _09862_ (.A1(_04857_),
    .A2(_04871_),
    .B1_N(_04858_),
    .X(_04935_));
 sky130_fd_sc_hd__xor2_4 _09863_ (.A(_04851_),
    .B(net89),
    .X(_04936_));
 sky130_fd_sc_hd__xor2_4 _09864_ (.A(_04935_),
    .B(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__or3_1 _09865_ (.A(_04856_),
    .B(_04934_),
    .C(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__nor2_1 _09866_ (.A(_04744_),
    .B(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand4_1 _09867_ (.A(net132),
    .B(_04597_),
    .C(_04646_),
    .D(_04649_),
    .Y(_04940_));
 sky130_fd_sc_hd__a31o_1 _09868_ (.A1(_04597_),
    .A2(_04646_),
    .A3(_04649_),
    .B1(net132),
    .X(_04941_));
 sky130_fd_sc_hd__nand3_1 _09869_ (.A(_04939_),
    .B(_04940_),
    .C(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__a21o_1 _09870_ (.A1(_04940_),
    .A2(_04941_),
    .B1(_04939_),
    .X(_04943_));
 sky130_fd_sc_hd__and3_1 _09871_ (.A(_04740_),
    .B(_04942_),
    .C(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__a21oi_1 _09872_ (.A1(_04942_),
    .A2(_04943_),
    .B1(_04740_),
    .Y(_04945_));
 sky130_fd_sc_hd__or3_1 _09873_ (.A(_04739_),
    .B(_04944_),
    .C(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__o21ai_1 _09874_ (.A1(_04944_),
    .A2(_04945_),
    .B1(_04739_),
    .Y(_04947_));
 sky130_fd_sc_hd__and3_1 _09875_ (.A(_04737_),
    .B(_04946_),
    .C(_04947_),
    .X(_04948_));
 sky130_fd_sc_hd__a21oi_1 _09876_ (.A1(_04946_),
    .A2(_04947_),
    .B1(_04737_),
    .Y(_04949_));
 sky130_fd_sc_hd__nor2_1 _09877_ (.A(_04728_),
    .B(_04733_),
    .Y(_04950_));
 sky130_fd_sc_hd__inv_2 _09878_ (.A(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__o211a_1 _09879_ (.A1(_04948_),
    .A2(_04949_),
    .B1(_04951_),
    .C1(_04735_),
    .X(_04952_));
 sky130_fd_sc_hd__a211o_1 _09880_ (.A1(_04951_),
    .A2(_04735_),
    .B1(_04948_),
    .C1(_04949_),
    .X(_04953_));
 sky130_fd_sc_hd__nand2_1 _09881_ (.A(_04463_),
    .B(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__inv_2 _09882_ (.A(\state[4] ),
    .Y(_04955_));
 sky130_fd_sc_hd__clkbuf_8 _09883_ (.A(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__nand2_1 _09884_ (.A(_04715_),
    .B(_04721_),
    .Y(_04957_));
 sky130_fd_sc_hd__or2b_1 _09885_ (.A(_04718_),
    .B_N(_04720_),
    .X(_04958_));
 sky130_fd_sc_hd__xor2_2 _09886_ (.A(net60),
    .B(net28),
    .X(_04959_));
 sky130_fd_sc_hd__xnor2_2 _09887_ (.A(net285),
    .B(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__xor2_1 _09888_ (.A(_04716_),
    .B(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__xnor2_1 _09889_ (.A(_04738_),
    .B(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__xnor2_1 _09890_ (.A(_04958_),
    .B(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__and3_1 _09891_ (.A(_04957_),
    .B(_04725_),
    .C(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__a21oi_1 _09892_ (.A1(_04957_),
    .A2(_04725_),
    .B1(_04963_),
    .Y(_04965_));
 sky130_fd_sc_hd__or3_1 _09893_ (.A(_04956_),
    .B(_04964_),
    .C(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__o21ai_4 _09894_ (.A1(_04952_),
    .A2(_04954_),
    .B1(_04966_),
    .Y(net167));
 sky130_fd_sc_hd__nand3_1 _09895_ (.A(_04737_),
    .B(_04946_),
    .C(_04947_),
    .Y(_04967_));
 sky130_fd_sc_hd__buf_2 _09896_ (.A(_04426_),
    .X(_04968_));
 sky130_fd_sc_hd__nor2_2 _09897_ (.A(_04739_),
    .B(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__and2_1 _09898_ (.A(_04739_),
    .B(_04968_),
    .X(_04970_));
 sky130_fd_sc_hd__or2_1 _09899_ (.A(_04969_),
    .B(_04970_),
    .X(_04971_));
 sky130_fd_sc_hd__clkbuf_2 _09900_ (.A(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__clkinv_8 _09901_ (.A(net133),
    .Y(_04973_));
 sky130_fd_sc_hd__a21bo_1 _09902_ (.A1(_04582_),
    .A2(_04646_),
    .B1_N(_04649_),
    .X(_04974_));
 sky130_fd_sc_hd__xnor2_2 _09903_ (.A(_04973_),
    .B(_04974_),
    .Y(_04975_));
 sky130_fd_sc_hd__or4_1 _09904_ (.A(_04910_),
    .B(_04856_),
    .C(_04934_),
    .D(_04937_),
    .X(_04976_));
 sky130_fd_sc_hd__nor2_2 _09905_ (.A(_04744_),
    .B(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__or4_1 _09906_ (.A(_04744_),
    .B(_04856_),
    .C(_04934_),
    .D(_04937_),
    .X(_04978_));
 sky130_fd_sc_hd__and2_1 _09907_ (.A(_04978_),
    .B(_04976_),
    .X(_04979_));
 sky130_fd_sc_hd__or2_1 _09908_ (.A(_04977_),
    .B(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__xor2_2 _09909_ (.A(_04975_),
    .B(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__and2_1 _09910_ (.A(_04940_),
    .B(_04942_),
    .X(_04982_));
 sky130_fd_sc_hd__xnor2_1 _09911_ (.A(_04981_),
    .B(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__xor2_1 _09912_ (.A(_04972_),
    .B(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__or2b_1 _09913_ (.A(_04944_),
    .B_N(_04946_),
    .X(_04985_));
 sky130_fd_sc_hd__xnor2_1 _09914_ (.A(_04984_),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__a21oi_2 _09915_ (.A1(_04967_),
    .A2(_04953_),
    .B1(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__a31o_1 _09916_ (.A1(_04967_),
    .A2(_04953_),
    .A3(_04986_),
    .B1(_04688_),
    .X(_04988_));
 sky130_fd_sc_hd__nor2_1 _09917_ (.A(_04958_),
    .B(_04962_),
    .Y(_04989_));
 sky130_fd_sc_hd__or2_1 _09918_ (.A(net61),
    .B(net29),
    .X(_04990_));
 sky130_fd_sc_hd__nand2_1 _09919_ (.A(net61),
    .B(net29),
    .Y(_04991_));
 sky130_fd_sc_hd__nand2_1 _09920_ (.A(_04990_),
    .B(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__nand2_1 _09921_ (.A(_04741_),
    .B(_04788_),
    .Y(_04993_));
 sky130_fd_sc_hd__or2_1 _09922_ (.A(_04741_),
    .B(_04788_),
    .X(_04994_));
 sky130_fd_sc_hd__and2_1 _09923_ (.A(_04993_),
    .B(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__xor2_1 _09924_ (.A(_04992_),
    .B(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__and2_1 _09925_ (.A(net60),
    .B(net28),
    .X(_04997_));
 sky130_fd_sc_hd__a21oi_2 _09926_ (.A1(net285),
    .A2(_04959_),
    .B1(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__xor2_1 _09927_ (.A(_04996_),
    .B(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__xnor2_1 _09928_ (.A(_04972_),
    .B(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__nor2_1 _09929_ (.A(_04716_),
    .B(_04960_),
    .Y(_05001_));
 sky130_fd_sc_hd__a21o_1 _09930_ (.A1(_04738_),
    .A2(_04961_),
    .B1(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__xnor2_1 _09931_ (.A(_05000_),
    .B(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__or3_1 _09932_ (.A(_04989_),
    .B(_04965_),
    .C(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__o21ai_1 _09933_ (.A1(_04989_),
    .A2(_04965_),
    .B1(_05003_),
    .Y(_05005_));
 sky130_fd_sc_hd__and2_1 _09934_ (.A(_05004_),
    .B(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__a2bb2o_4 _09935_ (.A1_N(_04987_),
    .A2_N(_04988_),
    .B1(_04444_),
    .B2(_05006_),
    .X(net168));
 sky130_fd_sc_hd__or2b_1 _09936_ (.A(_04982_),
    .B_N(_04981_),
    .X(_05007_));
 sky130_fd_sc_hd__nand2_1 _09937_ (.A(_04972_),
    .B(_04983_),
    .Y(_05008_));
 sky130_fd_sc_hd__and2_1 _09938_ (.A(_04738_),
    .B(_04968_),
    .X(_05009_));
 sky130_fd_sc_hd__clkbuf_4 _09939_ (.A(_04428_),
    .X(_05010_));
 sky130_fd_sc_hd__nand2_1 _09940_ (.A(_04968_),
    .B(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__or2_1 _09941_ (.A(_04968_),
    .B(_05010_),
    .X(_05012_));
 sky130_fd_sc_hd__and3_1 _09942_ (.A(_05009_),
    .B(_05011_),
    .C(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__a21oi_1 _09943_ (.A1(_05011_),
    .A2(_05012_),
    .B1(_05009_),
    .Y(_05014_));
 sky130_fd_sc_hd__nor2_2 _09944_ (.A(_05013_),
    .B(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__and3_1 _09945_ (.A(_04600_),
    .B(_04646_),
    .C(_04649_),
    .X(_05016_));
 sky130_fd_sc_hd__xnor2_1 _09946_ (.A(net134),
    .B(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__xnor2_4 _09947_ (.A(_04787_),
    .B(_04791_),
    .Y(_05018_));
 sky130_fd_sc_hd__or4_4 _09948_ (.A(_05018_),
    .B(_04856_),
    .C(_04934_),
    .D(_04937_),
    .X(_05019_));
 sky130_fd_sc_hd__nor2_2 _09949_ (.A(_04910_),
    .B(_05019_),
    .Y(_05020_));
 sky130_fd_sc_hd__or3_1 _09950_ (.A(_04912_),
    .B(_04938_),
    .C(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__mux2_1 _09951_ (.A0(_05021_),
    .A1(_05018_),
    .S(_04977_),
    .X(_05022_));
 sky130_fd_sc_hd__xor2_1 _09952_ (.A(_05017_),
    .B(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__o32a_1 _09953_ (.A1(_04975_),
    .A2(_04977_),
    .A3(_04979_),
    .B1(_04974_),
    .B2(_04973_),
    .X(_05024_));
 sky130_fd_sc_hd__xnor2_1 _09954_ (.A(_05023_),
    .B(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__xnor2_1 _09955_ (.A(_05015_),
    .B(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__nand3_1 _09956_ (.A(_05007_),
    .B(_05008_),
    .C(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__a21o_1 _09957_ (.A1(_05007_),
    .A2(_05008_),
    .B1(_05026_),
    .X(_05028_));
 sky130_fd_sc_hd__nand2_1 _09958_ (.A(_05027_),
    .B(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__and2_1 _09959_ (.A(_04984_),
    .B(_04985_),
    .X(_05030_));
 sky130_fd_sc_hd__or2_1 _09960_ (.A(_05030_),
    .B(_04987_),
    .X(_05031_));
 sky130_fd_sc_hd__xnor2_1 _09961_ (.A(_05029_),
    .B(_05031_),
    .Y(_05032_));
 sky130_fd_sc_hd__or2b_1 _09962_ (.A(_05000_),
    .B_N(_05002_),
    .X(_05033_));
 sky130_fd_sc_hd__or2_1 _09963_ (.A(net62),
    .B(net30),
    .X(_05034_));
 sky130_fd_sc_hd__nand2_1 _09964_ (.A(net62),
    .B(net30),
    .Y(_05035_));
 sky130_fd_sc_hd__nand2_1 _09965_ (.A(_05034_),
    .B(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__xor2_1 _09966_ (.A(_04784_),
    .B(_04788_),
    .X(_05037_));
 sky130_fd_sc_hd__mux2_1 _09967_ (.A0(_04784_),
    .A1(_05037_),
    .S(_04993_),
    .X(_05038_));
 sky130_fd_sc_hd__xor2_1 _09968_ (.A(_05036_),
    .B(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__a21boi_1 _09969_ (.A1(_04990_),
    .A2(_04995_),
    .B1_N(_04991_),
    .Y(_05040_));
 sky130_fd_sc_hd__nor2_1 _09970_ (.A(_05039_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__and2_1 _09971_ (.A(_05039_),
    .B(_05040_),
    .X(_05042_));
 sky130_fd_sc_hd__nor2_1 _09972_ (.A(_05041_),
    .B(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__xnor2_1 _09973_ (.A(_05015_),
    .B(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__nor2_1 _09974_ (.A(_04996_),
    .B(_04998_),
    .Y(_05045_));
 sky130_fd_sc_hd__a21o_1 _09975_ (.A1(_04972_),
    .A2(_04999_),
    .B1(_05045_),
    .X(_05046_));
 sky130_fd_sc_hd__xor2_1 _09976_ (.A(_05044_),
    .B(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__and3_1 _09977_ (.A(_05033_),
    .B(_05005_),
    .C(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__a21oi_1 _09978_ (.A1(_05033_),
    .A2(_05005_),
    .B1(_05047_),
    .Y(_05049_));
 sky130_fd_sc_hd__nor2_1 _09979_ (.A(_05048_),
    .B(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__a22o_4 _09980_ (.A1(_04464_),
    .A2(_05032_),
    .B1(_05050_),
    .B2(_04444_),
    .X(net169));
 sky130_fd_sc_hd__buf_2 _09981_ (.A(\pixel_cnt[7] ),
    .X(_05051_));
 sky130_fd_sc_hd__buf_2 _09982_ (.A(\pixel_cnt[6] ),
    .X(_05052_));
 sky130_fd_sc_hd__buf_2 _09983_ (.A(\pixel_cnt[4] ),
    .X(_05053_));
 sky130_fd_sc_hd__buf_2 _09984_ (.A(\pixel_cnt[5] ),
    .X(_05054_));
 sky130_fd_sc_hd__and4bb_4 _09985_ (.A_N(_05051_),
    .B_N(_05052_),
    .C(_05053_),
    .D(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__clkbuf_8 _09986_ (.A(_05055_),
    .X(_05056_));
 sky130_fd_sc_hd__buf_6 _09987_ (.A(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__buf_8 _09988_ (.A(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__buf_6 _09989_ (.A(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__or2b_1 _09990_ (.A(_04968_),
    .B_N(_05010_),
    .X(_05060_));
 sky130_fd_sc_hd__clkbuf_4 _09991_ (.A(_04427_),
    .X(_05061_));
 sky130_fd_sc_hd__nand2_1 _09992_ (.A(_04738_),
    .B(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__or2_1 _09993_ (.A(_04738_),
    .B(_05061_),
    .X(_05063_));
 sky130_fd_sc_hd__a21oi_1 _09994_ (.A1(_05062_),
    .A2(_05063_),
    .B1(_05060_),
    .Y(_05064_));
 sky130_fd_sc_hd__a311o_1 _09995_ (.A1(_05060_),
    .A2(_05062_),
    .A3(_05063_),
    .B1(_05064_),
    .C1(_05013_),
    .X(_05065_));
 sky130_fd_sc_hd__nand2b_2 _09996_ (.A_N(_05059_),
    .B(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__inv_2 _09997_ (.A(net135),
    .Y(_05067_));
 sky130_fd_sc_hd__a21bo_1 _09998_ (.A1(_04580_),
    .A2(_04646_),
    .B1_N(_04649_),
    .X(_05068_));
 sky130_fd_sc_hd__xnor2_1 _09999_ (.A(_05067_),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__a21oi_1 _10000_ (.A1(_05018_),
    .A2(_04977_),
    .B1(_05020_),
    .Y(_05070_));
 sky130_fd_sc_hd__inv_2 _10001_ (.A(_04744_),
    .Y(_05071_));
 sky130_fd_sc_hd__mux2_2 _10002_ (.A0(_05071_),
    .A1(_04978_),
    .S(_05019_),
    .X(_05072_));
 sky130_fd_sc_hd__nor2_1 _10003_ (.A(_04915_),
    .B(_04938_),
    .Y(_05073_));
 sky130_fd_sc_hd__xnor2_2 _10004_ (.A(_05072_),
    .B(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__and2b_1 _10005_ (.A_N(_05070_),
    .B(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__and2b_1 _10006_ (.A_N(_05074_),
    .B(_05070_),
    .X(_05076_));
 sky130_fd_sc_hd__nor2_1 _10007_ (.A(_05075_),
    .B(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__xnor2_1 _10008_ (.A(_05069_),
    .B(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__nor2_1 _10009_ (.A(_05017_),
    .B(_05022_),
    .Y(_05079_));
 sky130_fd_sc_hd__a21o_1 _10010_ (.A1(net134),
    .A2(_05016_),
    .B1(_05079_),
    .X(_05080_));
 sky130_fd_sc_hd__xor2_1 _10011_ (.A(_05078_),
    .B(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__xor2_1 _10012_ (.A(_05066_),
    .B(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__and2_1 _10013_ (.A(_05017_),
    .B(_05022_),
    .X(_05083_));
 sky130_fd_sc_hd__nand2_1 _10014_ (.A(_05015_),
    .B(_05025_),
    .Y(_05084_));
 sky130_fd_sc_hd__o31a_1 _10015_ (.A1(_05083_),
    .A2(_05079_),
    .A3(_05024_),
    .B1(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__xor2_1 _10016_ (.A(_05082_),
    .B(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__inv_2 _10017_ (.A(_05028_),
    .Y(_05087_));
 sky130_fd_sc_hd__o21a_1 _10018_ (.A1(_05087_),
    .A2(_05031_),
    .B1(_05027_),
    .X(_05088_));
 sky130_fd_sc_hd__o21ai_1 _10019_ (.A1(_05086_),
    .A2(_05088_),
    .B1(_04464_),
    .Y(_05089_));
 sky130_fd_sc_hd__o311a_2 _10020_ (.A1(_05030_),
    .A2(_04987_),
    .A3(_05087_),
    .B1(_05086_),
    .C1(_05027_),
    .X(_05090_));
 sky130_fd_sc_hd__and2b_1 _10021_ (.A_N(_05044_),
    .B(_05046_),
    .X(_05091_));
 sky130_fd_sc_hd__or2_1 _10022_ (.A(net63),
    .B(net31),
    .X(_05092_));
 sky130_fd_sc_hd__nand2_1 _10023_ (.A(net63),
    .B(net31),
    .Y(_05093_));
 sky130_fd_sc_hd__nand2_1 _10024_ (.A(_05092_),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__xor2_2 _10025_ (.A(_04741_),
    .B(net90),
    .X(_05095_));
 sky130_fd_sc_hd__o21ai_2 _10026_ (.A1(_04741_),
    .A2(_04784_),
    .B1(_05037_),
    .Y(_05096_));
 sky130_fd_sc_hd__xnor2_2 _10027_ (.A(_05095_),
    .B(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__xor2_1 _10028_ (.A(_05094_),
    .B(_05097_),
    .X(_05098_));
 sky130_fd_sc_hd__a21bo_1 _10029_ (.A1(_05034_),
    .A2(_05038_),
    .B1_N(_05035_),
    .X(_05099_));
 sky130_fd_sc_hd__and2b_1 _10030_ (.A_N(_05098_),
    .B(_05099_),
    .X(_05100_));
 sky130_fd_sc_hd__and2b_1 _10031_ (.A_N(_05099_),
    .B(_05098_),
    .X(_05101_));
 sky130_fd_sc_hd__nor2_1 _10032_ (.A(_05100_),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__xor2_1 _10033_ (.A(_05066_),
    .B(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__a21o_1 _10034_ (.A1(_05015_),
    .A2(_05043_),
    .B1(_05041_),
    .X(_05104_));
 sky130_fd_sc_hd__xnor2_1 _10035_ (.A(_05103_),
    .B(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__o21a_1 _10036_ (.A1(_05091_),
    .A2(_05049_),
    .B1(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__nor2_1 _10037_ (.A(_04956_),
    .B(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__or3_1 _10038_ (.A(_05091_),
    .B(_05049_),
    .C(_05105_),
    .X(_05108_));
 sky130_fd_sc_hd__a2bb2o_4 _10039_ (.A1_N(_05089_),
    .A2_N(_05090_),
    .B1(_05107_),
    .B2(_05108_),
    .X(net170));
 sky130_fd_sc_hd__nor2_1 _10040_ (.A(_05082_),
    .B(_05085_),
    .Y(_05109_));
 sky130_fd_sc_hd__and2b_1 _10041_ (.A_N(_05010_),
    .B(_05061_),
    .X(_05110_));
 sky130_fd_sc_hd__or2_2 _10042_ (.A(_04969_),
    .B(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__and2b_1 _10043_ (.A_N(_05061_),
    .B(_05010_),
    .X(_05112_));
 sky130_fd_sc_hd__o21ba_1 _10044_ (.A1(_04969_),
    .A2(_04970_),
    .B1_N(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__xnor2_4 _10045_ (.A(_05111_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__nand2_1 _10046_ (.A(_05020_),
    .B(_05074_),
    .Y(_05115_));
 sky130_fd_sc_hd__or4_2 _10047_ (.A(_04915_),
    .B(_04856_),
    .C(_04934_),
    .D(_04937_),
    .X(_05116_));
 sky130_fd_sc_hd__o22ai_4 _10048_ (.A1(_04744_),
    .A2(_05019_),
    .B1(_05072_),
    .B2(net287),
    .Y(_05117_));
 sky130_fd_sc_hd__mux2_2 _10049_ (.A0(_04911_),
    .A1(_04976_),
    .S(_05116_),
    .X(_05118_));
 sky130_fd_sc_hd__or4_1 _10050_ (.A(_04906_),
    .B(_04856_),
    .C(_04934_),
    .D(_04937_),
    .X(_05119_));
 sky130_fd_sc_hd__buf_6 _10051_ (.A(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__xnor2_2 _10052_ (.A(_05118_),
    .B(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__xnor2_2 _10053_ (.A(_05117_),
    .B(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__xor2_1 _10054_ (.A(_05115_),
    .B(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__and3_1 _10055_ (.A(_05018_),
    .B(_04977_),
    .C(_05074_),
    .X(_05124_));
 sky130_fd_sc_hd__xnor2_2 _10056_ (.A(_05123_),
    .B(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__xnor2_2 _10057_ (.A(net136),
    .B(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__o32a_1 _10058_ (.A1(_05069_),
    .A2(_05075_),
    .A3(_05076_),
    .B1(_05068_),
    .B2(_05067_),
    .X(_05127_));
 sky130_fd_sc_hd__xnor2_1 _10059_ (.A(_05126_),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__xnor2_1 _10060_ (.A(_05114_),
    .B(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__and2b_1 _10061_ (.A_N(_05066_),
    .B(_05081_),
    .X(_05130_));
 sky130_fd_sc_hd__a21o_1 _10062_ (.A1(_05078_),
    .A2(_05080_),
    .B1(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__and2b_1 _10063_ (.A_N(_05129_),
    .B(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__or2b_1 _10064_ (.A(_05131_),
    .B_N(_05129_),
    .X(_05133_));
 sky130_fd_sc_hd__and2b_1 _10065_ (.A_N(_05132_),
    .B(_05133_),
    .X(_05134_));
 sky130_fd_sc_hd__or3_1 _10066_ (.A(_05109_),
    .B(_05090_),
    .C(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__o21ai_1 _10067_ (.A1(_05109_),
    .A2(_05090_),
    .B1(_05134_),
    .Y(_05136_));
 sky130_fd_sc_hd__and2b_1 _10068_ (.A_N(_05103_),
    .B(_05104_),
    .X(_05137_));
 sky130_fd_sc_hd__and2b_1 _10069_ (.A_N(_05066_),
    .B(_05102_),
    .X(_05138_));
 sky130_fd_sc_hd__or2_1 _10070_ (.A(net64),
    .B(net32),
    .X(_05139_));
 sky130_fd_sc_hd__nand2_1 _10071_ (.A(net64),
    .B(net32),
    .Y(_05140_));
 sky130_fd_sc_hd__nand2_1 _10072_ (.A(_05139_),
    .B(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand2_2 _10073_ (.A(_04784_),
    .B(_05095_),
    .Y(_05142_));
 sky130_fd_sc_hd__or2b_1 _10074_ (.A(_04741_),
    .B_N(net90),
    .X(_05143_));
 sky130_fd_sc_hd__xor2_2 _10075_ (.A(net91),
    .B(_04788_),
    .X(_05144_));
 sky130_fd_sc_hd__xnor2_2 _10076_ (.A(_05143_),
    .B(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__xnor2_4 _10077_ (.A(_05142_),
    .B(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__nand2_1 _10078_ (.A(_04784_),
    .B(_04788_),
    .Y(_05147_));
 sky130_fd_sc_hd__o32a_2 _10079_ (.A1(net90),
    .A2(_04784_),
    .A3(_04993_),
    .B1(_05147_),
    .B2(_05095_),
    .X(_05148_));
 sky130_fd_sc_hd__xnor2_4 _10080_ (.A(_05146_),
    .B(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__xor2_2 _10081_ (.A(_05141_),
    .B(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__a21bo_1 _10082_ (.A1(_05092_),
    .A2(_05097_),
    .B1_N(_05093_),
    .X(_05151_));
 sky130_fd_sc_hd__xnor2_2 _10083_ (.A(_05150_),
    .B(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__xnor2_1 _10084_ (.A(_05114_),
    .B(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__o21ai_1 _10085_ (.A1(_05100_),
    .A2(_05138_),
    .B1(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__or3_1 _10086_ (.A(_05100_),
    .B(_05138_),
    .C(_05153_),
    .X(_05155_));
 sky130_fd_sc_hd__and2_1 _10087_ (.A(_05154_),
    .B(_05155_),
    .X(_05156_));
 sky130_fd_sc_hd__or3_1 _10088_ (.A(_05137_),
    .B(_05106_),
    .C(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__o21ai_1 _10089_ (.A1(_05137_),
    .A2(_05106_),
    .B1(_05156_),
    .Y(_05158_));
 sky130_fd_sc_hd__and3_1 _10090_ (.A(_04443_),
    .B(_05157_),
    .C(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__a31o_2 _10091_ (.A1(_04464_),
    .A2(_05135_),
    .A3(_05136_),
    .B1(_05159_),
    .X(net171));
 sky130_fd_sc_hd__nand2_1 _10092_ (.A(_04738_),
    .B(_04968_),
    .Y(_05160_));
 sky130_fd_sc_hd__o21ai_1 _10093_ (.A1(_04738_),
    .A2(_04968_),
    .B1(_05110_),
    .Y(_05161_));
 sky130_fd_sc_hd__o221a_2 _10094_ (.A1(_05061_),
    .A2(_05060_),
    .B1(_05112_),
    .B2(_05160_),
    .C1(_05161_),
    .X(_05162_));
 sky130_fd_sc_hd__nand2_1 _10095_ (.A(net136),
    .B(_05125_),
    .Y(_05163_));
 sky130_fd_sc_hd__and4_1 _10096_ (.A(_05018_),
    .B(_04977_),
    .C(_05074_),
    .D(_05122_),
    .X(_05164_));
 sky130_fd_sc_hd__a31o_1 _10097_ (.A1(_05020_),
    .A2(_05074_),
    .A3(_05122_),
    .B1(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__and2b_1 _10098_ (.A_N(_05121_),
    .B(_05117_),
    .X(_05166_));
 sky130_fd_sc_hd__mux2_1 _10099_ (.A0(_04907_),
    .A1(_05019_),
    .S(_05120_),
    .X(_05167_));
 sky130_fd_sc_hd__xnor2_1 _10100_ (.A(_04935_),
    .B(_04936_),
    .Y(_05168_));
 sky130_fd_sc_hd__o31a_1 _10101_ (.A1(_04903_),
    .A2(_04856_),
    .A3(_04934_),
    .B1(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__xnor2_1 _10102_ (.A(_05167_),
    .B(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__o22ai_2 _10103_ (.A1(_04910_),
    .A2(net287),
    .B1(_05118_),
    .B2(_05120_),
    .Y(_05171_));
 sky130_fd_sc_hd__xor2_1 _10104_ (.A(_05170_),
    .B(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__or2_1 _10105_ (.A(_05166_),
    .B(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__nand2_1 _10106_ (.A(_05166_),
    .B(_05172_),
    .Y(_05174_));
 sky130_fd_sc_hd__nand2_1 _10107_ (.A(_05173_),
    .B(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__xnor2_1 _10108_ (.A(_05165_),
    .B(_05175_),
    .Y(_05176_));
 sky130_fd_sc_hd__xnor2_1 _10109_ (.A(net106),
    .B(_05176_),
    .Y(_05177_));
 sky130_fd_sc_hd__xnor2_1 _10110_ (.A(_05163_),
    .B(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__xor2_1 _10111_ (.A(_05162_),
    .B(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__o22ai_2 _10112_ (.A1(_05126_),
    .A2(_05127_),
    .B1(_05128_),
    .B2(_05114_),
    .Y(_05180_));
 sky130_fd_sc_hd__xnor2_1 _10113_ (.A(_05179_),
    .B(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__o31ai_2 _10114_ (.A1(_05109_),
    .A2(_05090_),
    .A3(_05132_),
    .B1(_05133_),
    .Y(_05182_));
 sky130_fd_sc_hd__nor2_1 _10115_ (.A(_05181_),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__a21o_1 _10116_ (.A1(_05181_),
    .A2(_05182_),
    .B1(_04688_),
    .X(_05184_));
 sky130_fd_sc_hd__or2_1 _10117_ (.A(net34),
    .B(net2),
    .X(_05185_));
 sky130_fd_sc_hd__nand2_1 _10118_ (.A(net34),
    .B(net2),
    .Y(_05186_));
 sky130_fd_sc_hd__nand2_1 _10119_ (.A(_05185_),
    .B(_05186_),
    .Y(_05187_));
 sky130_fd_sc_hd__or2b_1 _10120_ (.A(_05142_),
    .B_N(_05145_),
    .X(_05188_));
 sky130_fd_sc_hd__or2b_1 _10121_ (.A(_05148_),
    .B_N(_05146_),
    .X(_05189_));
 sky130_fd_sc_hd__o21a_1 _10122_ (.A1(_04741_),
    .A2(_05144_),
    .B1(net90),
    .X(_05190_));
 sky130_fd_sc_hd__xor2_1 _10123_ (.A(net92),
    .B(_04784_),
    .X(_05191_));
 sky130_fd_sc_hd__nor2_1 _10124_ (.A(_04788_),
    .B(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__inv_2 _10125_ (.A(net91),
    .Y(_05193_));
 sky130_fd_sc_hd__o21a_1 _10126_ (.A1(_05193_),
    .A2(_04788_),
    .B1(_05191_),
    .X(_05194_));
 sky130_fd_sc_hd__a21oi_1 _10127_ (.A1(net91),
    .A2(_05192_),
    .B1(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__xor2_1 _10128_ (.A(_05190_),
    .B(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__a21o_1 _10129_ (.A1(_05188_),
    .A2(_05189_),
    .B1(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__nand3_1 _10130_ (.A(_05188_),
    .B(_05189_),
    .C(_05196_),
    .Y(_05198_));
 sky130_fd_sc_hd__and2_2 _10131_ (.A(_05197_),
    .B(_05198_),
    .X(_05199_));
 sky130_fd_sc_hd__xor2_1 _10132_ (.A(_05187_),
    .B(_05199_),
    .X(_05200_));
 sky130_fd_sc_hd__a21boi_1 _10133_ (.A1(_05139_),
    .A2(_05149_),
    .B1_N(_05140_),
    .Y(_05201_));
 sky130_fd_sc_hd__xnor2_1 _10134_ (.A(_05200_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__xnor2_1 _10135_ (.A(_05202_),
    .B(_05162_),
    .Y(_05203_));
 sky130_fd_sc_hd__inv_2 _10136_ (.A(_05151_),
    .Y(_05204_));
 sky130_fd_sc_hd__inv_2 _10137_ (.A(_05152_),
    .Y(_05205_));
 sky130_fd_sc_hd__o22a_1 _10138_ (.A1(_05150_),
    .A2(_05204_),
    .B1(_05205_),
    .B2(_05114_),
    .X(_05206_));
 sky130_fd_sc_hd__xnor2_1 _10139_ (.A(_05203_),
    .B(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__and3_1 _10140_ (.A(_05154_),
    .B(_05158_),
    .C(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__a21oi_1 _10141_ (.A1(_05154_),
    .A2(_05158_),
    .B1(_05207_),
    .Y(_05209_));
 sky130_fd_sc_hd__or3_1 _10142_ (.A(_04956_),
    .B(_05208_),
    .C(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__o21ai_4 _10143_ (.A1(_05183_),
    .A2(_05184_),
    .B1(_05210_),
    .Y(net141));
 sky130_fd_sc_hd__nand2_1 _10144_ (.A(_05179_),
    .B(_05180_),
    .Y(_05211_));
 sky130_fd_sc_hd__inv_2 _10145_ (.A(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__nand2_2 _10146_ (.A(_05061_),
    .B(_05010_),
    .Y(_05213_));
 sky130_fd_sc_hd__a21o_1 _10147_ (.A1(_04968_),
    .A2(_05010_),
    .B1(_05061_),
    .X(_05214_));
 sky130_fd_sc_hd__nand2_2 _10148_ (.A(_05213_),
    .B(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__nand2_1 _10149_ (.A(net106),
    .B(_05176_),
    .Y(_05216_));
 sky130_fd_sc_hd__nand2_1 _10150_ (.A(_05170_),
    .B(_05171_),
    .Y(_05217_));
 sky130_fd_sc_hd__nand2_1 _10151_ (.A(_05019_),
    .B(_05120_),
    .Y(_05218_));
 sky130_fd_sc_hd__o2bb2a_1 _10152_ (.A1_N(_05218_),
    .A2_N(_05169_),
    .B1(_05018_),
    .B2(_05120_),
    .X(_05219_));
 sky130_fd_sc_hd__mux2_1 _10153_ (.A0(_04904_),
    .A1(_05169_),
    .S(_05116_),
    .X(_05220_));
 sky130_fd_sc_hd__nor2_2 _10154_ (.A(_04856_),
    .B(net283),
    .Y(_05221_));
 sky130_fd_sc_hd__a21oi_2 _10155_ (.A1(_04901_),
    .A2(_05221_),
    .B1(_04937_),
    .Y(_05222_));
 sky130_fd_sc_hd__xnor2_1 _10156_ (.A(_05220_),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__xnor2_1 _10157_ (.A(_05219_),
    .B(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__nor2_1 _10158_ (.A(_05217_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__and2_1 _10159_ (.A(_05217_),
    .B(_05224_),
    .X(_05226_));
 sky130_fd_sc_hd__nor2_1 _10160_ (.A(_05225_),
    .B(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__a31o_1 _10161_ (.A1(_05020_),
    .A2(_05074_),
    .A3(_05122_),
    .B1(_05166_),
    .X(_05228_));
 sky130_fd_sc_hd__a22o_1 _10162_ (.A1(_05164_),
    .A2(_05173_),
    .B1(_05228_),
    .B2(_05172_),
    .X(_05229_));
 sky130_fd_sc_hd__xor2_1 _10163_ (.A(_05227_),
    .B(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__xnor2_1 _10164_ (.A(net107),
    .B(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__xnor2_1 _10165_ (.A(_05216_),
    .B(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__xnor2_1 _10166_ (.A(_05215_),
    .B(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__or2_1 _10167_ (.A(_05163_),
    .B(_05177_),
    .X(_05234_));
 sky130_fd_sc_hd__o21ai_1 _10168_ (.A1(_05162_),
    .A2(_05178_),
    .B1(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__xnor2_1 _10169_ (.A(_05233_),
    .B(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__or3_1 _10170_ (.A(_05212_),
    .B(_05183_),
    .C(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__o21ai_1 _10171_ (.A1(_05212_),
    .A2(_05183_),
    .B1(_05236_),
    .Y(_05238_));
 sky130_fd_sc_hd__nor2_1 _10172_ (.A(_05203_),
    .B(_05206_),
    .Y(_05239_));
 sky130_fd_sc_hd__or2_1 _10173_ (.A(net35),
    .B(net3),
    .X(_05240_));
 sky130_fd_sc_hd__nand2_1 _10174_ (.A(net35),
    .B(net3),
    .Y(_05241_));
 sky130_fd_sc_hd__nand2_1 _10175_ (.A(_05240_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__or2b_1 _10176_ (.A(_05195_),
    .B_N(_05190_),
    .X(_05243_));
 sky130_fd_sc_hd__or2_1 _10177_ (.A(_05193_),
    .B(_05192_),
    .X(_05244_));
 sky130_fd_sc_hd__xor2_1 _10178_ (.A(_04781_),
    .B(net90),
    .X(_05245_));
 sky130_fd_sc_hd__nor2_1 _10179_ (.A(_04784_),
    .B(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__inv_2 _10180_ (.A(net92),
    .Y(_05247_));
 sky130_fd_sc_hd__o21a_1 _10181_ (.A1(_05247_),
    .A2(_04784_),
    .B1(_05245_),
    .X(_05248_));
 sky130_fd_sc_hd__a21oi_1 _10182_ (.A1(net92),
    .A2(_05246_),
    .B1(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__or2_1 _10183_ (.A(_05244_),
    .B(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__nand2_1 _10184_ (.A(_05244_),
    .B(_05249_),
    .Y(_05251_));
 sky130_fd_sc_hd__nand2_1 _10185_ (.A(_05250_),
    .B(_05251_),
    .Y(_05252_));
 sky130_fd_sc_hd__a21o_1 _10186_ (.A1(_05243_),
    .A2(_05197_),
    .B1(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__nand3_1 _10187_ (.A(_05243_),
    .B(_05197_),
    .C(_05252_),
    .Y(_05254_));
 sky130_fd_sc_hd__and2_2 _10188_ (.A(_05253_),
    .B(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__xor2_1 _10189_ (.A(_05242_),
    .B(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__a21boi_1 _10190_ (.A1(_05185_),
    .A2(_05199_),
    .B1_N(_05186_),
    .Y(_05257_));
 sky130_fd_sc_hd__xor2_1 _10191_ (.A(_05256_),
    .B(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__xnor2_1 _10192_ (.A(_05215_),
    .B(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__or2_1 _10193_ (.A(_05200_),
    .B(_05201_),
    .X(_05260_));
 sky130_fd_sc_hd__o21a_1 _10194_ (.A1(_05202_),
    .A2(_05162_),
    .B1(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__xnor2_1 _10195_ (.A(_05259_),
    .B(_05261_),
    .Y(_05262_));
 sky130_fd_sc_hd__or3_1 _10196_ (.A(_05239_),
    .B(_05209_),
    .C(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__o21ai_1 _10197_ (.A1(_05239_),
    .A2(_05209_),
    .B1(_05262_),
    .Y(_05264_));
 sky130_fd_sc_hd__and3_1 _10198_ (.A(_04443_),
    .B(_05263_),
    .C(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__a31o_4 _10199_ (.A1(_04464_),
    .A2(_05237_),
    .A3(_05238_),
    .B1(_05265_),
    .X(net142));
 sky130_fd_sc_hd__or2b_1 _10200_ (.A(_05261_),
    .B_N(_05259_),
    .X(_05266_));
 sky130_fd_sc_hd__or2_1 _10201_ (.A(net36),
    .B(net4),
    .X(_05267_));
 sky130_fd_sc_hd__nand2_1 _10202_ (.A(net36),
    .B(net4),
    .Y(_05268_));
 sky130_fd_sc_hd__nand2_1 _10203_ (.A(_05267_),
    .B(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__xor2_1 _10204_ (.A(_04780_),
    .B(net91),
    .X(_05270_));
 sky130_fd_sc_hd__nor2_1 _10205_ (.A(net90),
    .B(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__inv_2 _10206_ (.A(net284),
    .Y(_05272_));
 sky130_fd_sc_hd__o21a_1 _10207_ (.A1(_05272_),
    .A2(net90),
    .B1(_05270_),
    .X(_05273_));
 sky130_fd_sc_hd__a21oi_1 _10208_ (.A1(net284),
    .A2(_05271_),
    .B1(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__or3_1 _10209_ (.A(_05247_),
    .B(_05246_),
    .C(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__o21ai_1 _10210_ (.A1(_05247_),
    .A2(_05246_),
    .B1(_05274_),
    .Y(_05276_));
 sky130_fd_sc_hd__nand2_1 _10211_ (.A(_05275_),
    .B(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hd__a21o_1 _10212_ (.A1(_05250_),
    .A2(_05253_),
    .B1(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__nand3_1 _10213_ (.A(_05250_),
    .B(_05253_),
    .C(_05277_),
    .Y(_05279_));
 sky130_fd_sc_hd__and2_2 _10214_ (.A(_05278_),
    .B(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__xor2_1 _10215_ (.A(_05269_),
    .B(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__a21boi_1 _10216_ (.A1(_05240_),
    .A2(_05255_),
    .B1_N(_05241_),
    .Y(_05282_));
 sky130_fd_sc_hd__xor2_1 _10217_ (.A(_05281_),
    .B(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__xnor2_1 _10218_ (.A(_05213_),
    .B(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__nor2_1 _10219_ (.A(_05256_),
    .B(_05257_),
    .Y(_05285_));
 sky130_fd_sc_hd__a31o_1 _10220_ (.A1(_05213_),
    .A2(_05214_),
    .A3(_05258_),
    .B1(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__xnor2_1 _10221_ (.A(_05284_),
    .B(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__and3_1 _10222_ (.A(_05266_),
    .B(_05264_),
    .C(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__a21o_1 _10223_ (.A1(_05266_),
    .A2(_05264_),
    .B1(_05287_),
    .X(_05289_));
 sky130_fd_sc_hd__nand2_1 _10224_ (.A(_04724_),
    .B(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__or3b_1 _10225_ (.A(_05181_),
    .B(_05182_),
    .C_N(_05236_),
    .X(_05291_));
 sky130_fd_sc_hd__and2b_1 _10226_ (.A_N(_05235_),
    .B(net281),
    .X(_05292_));
 sky130_fd_sc_hd__or2b_1 _10227_ (.A(net281),
    .B_N(_05235_),
    .X(_05293_));
 sky130_fd_sc_hd__o21a_1 _10228_ (.A1(_05211_),
    .A2(_05292_),
    .B1(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__nand2_1 _10229_ (.A(net107),
    .B(_05230_),
    .Y(_05295_));
 sky130_fd_sc_hd__a21oi_1 _10230_ (.A1(_05227_),
    .A2(_05229_),
    .B1(_05225_),
    .Y(_05296_));
 sky130_fd_sc_hd__nor2_1 _10231_ (.A(_05219_),
    .B(_05223_),
    .Y(_05297_));
 sky130_fd_sc_hd__mux2_1 _10232_ (.A0(_04901_),
    .A1(_05222_),
    .S(_05120_),
    .X(_05298_));
 sky130_fd_sc_hd__a21oi_4 _10233_ (.A1(_04899_),
    .A2(_05221_),
    .B1(_04937_),
    .Y(_05299_));
 sky130_fd_sc_hd__xnor2_2 _10234_ (.A(_05298_),
    .B(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__a22o_1 _10235_ (.A1(_04903_),
    .A2(_05073_),
    .B1(_05220_),
    .B2(_05222_),
    .X(_05301_));
 sky130_fd_sc_hd__xnor2_2 _10236_ (.A(_05300_),
    .B(_05301_),
    .Y(_05302_));
 sky130_fd_sc_hd__xor2_2 _10237_ (.A(_05297_),
    .B(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__xnor2_1 _10238_ (.A(_05296_),
    .B(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__xnor2_1 _10239_ (.A(net108),
    .B(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__xor2_1 _10240_ (.A(_05295_),
    .B(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__xnor2_1 _10241_ (.A(_05213_),
    .B(_05306_),
    .Y(_05307_));
 sky130_fd_sc_hd__or2_1 _10242_ (.A(_05216_),
    .B(_05231_),
    .X(_05308_));
 sky130_fd_sc_hd__o21ai_1 _10243_ (.A1(_05215_),
    .A2(_05232_),
    .B1(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__xnor2_1 _10244_ (.A(_05307_),
    .B(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__a21o_1 _10245_ (.A1(_05291_),
    .A2(_05294_),
    .B1(_05310_),
    .X(_05311_));
 sky130_fd_sc_hd__nand2_1 _10246_ (.A(_04463_),
    .B(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__a31o_1 _10247_ (.A1(_05291_),
    .A2(_05294_),
    .A3(_05310_),
    .B1(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__o21ai_4 _10248_ (.A1(_05288_),
    .A2(_05290_),
    .B1(_05313_),
    .Y(net143));
 sky130_fd_sc_hd__nand2_1 _10249_ (.A(_05284_),
    .B(_05286_),
    .Y(_05314_));
 sky130_fd_sc_hd__or2_1 _10250_ (.A(net37),
    .B(net5),
    .X(_05315_));
 sky130_fd_sc_hd__nand2_1 _10251_ (.A(net37),
    .B(net5),
    .Y(_05316_));
 sky130_fd_sc_hd__nand2_1 _10252_ (.A(_05315_),
    .B(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__xor2_1 _10253_ (.A(_04807_),
    .B(net92),
    .X(_05318_));
 sky130_fd_sc_hd__nor2_1 _10254_ (.A(net91),
    .B(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hd__inv_2 _10255_ (.A(_04780_),
    .Y(_05320_));
 sky130_fd_sc_hd__o21a_1 _10256_ (.A1(_05320_),
    .A2(net91),
    .B1(_05318_),
    .X(_05321_));
 sky130_fd_sc_hd__a21oi_1 _10257_ (.A1(_04780_),
    .A2(_05319_),
    .B1(_05321_),
    .Y(_05322_));
 sky130_fd_sc_hd__or3_1 _10258_ (.A(_05272_),
    .B(_05271_),
    .C(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__o21ai_1 _10259_ (.A1(_05272_),
    .A2(_05271_),
    .B1(_05322_),
    .Y(_05324_));
 sky130_fd_sc_hd__nand2_1 _10260_ (.A(_05323_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__a21o_1 _10261_ (.A1(_05275_),
    .A2(_05278_),
    .B1(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__nand3_1 _10262_ (.A(_05275_),
    .B(_05278_),
    .C(_05325_),
    .Y(_05327_));
 sky130_fd_sc_hd__and2_2 _10263_ (.A(_05326_),
    .B(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__xor2_1 _10264_ (.A(_05317_),
    .B(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__a21boi_1 _10265_ (.A1(_05267_),
    .A2(_05280_),
    .B1_N(_05268_),
    .Y(_05330_));
 sky130_fd_sc_hd__nor2_1 _10266_ (.A(_05329_),
    .B(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__and2_1 _10267_ (.A(_05329_),
    .B(_05330_),
    .X(_05332_));
 sky130_fd_sc_hd__nor2_1 _10268_ (.A(_05331_),
    .B(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__and3_1 _10269_ (.A(_05061_),
    .B(_05010_),
    .C(_05283_),
    .X(_05334_));
 sky130_fd_sc_hd__o21ba_1 _10270_ (.A1(_05281_),
    .A2(_05282_),
    .B1_N(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__xor2_1 _10271_ (.A(_05333_),
    .B(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__and3_1 _10272_ (.A(_05314_),
    .B(_05289_),
    .C(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__a21o_1 _10273_ (.A1(_05314_),
    .A2(_05289_),
    .B1(_05336_),
    .X(_05338_));
 sky130_fd_sc_hd__nand2_1 _10274_ (.A(_04724_),
    .B(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__nand2_1 _10275_ (.A(_05307_),
    .B(_05309_),
    .Y(_05340_));
 sky130_fd_sc_hd__nor2_1 _10276_ (.A(_05295_),
    .B(_05305_),
    .Y(_05341_));
 sky130_fd_sc_hd__and3_1 _10277_ (.A(_05061_),
    .B(_05010_),
    .C(_05306_),
    .X(_05342_));
 sky130_fd_sc_hd__nand2_1 _10278_ (.A(net108),
    .B(_05304_),
    .Y(_05343_));
 sky130_fd_sc_hd__or2b_1 _10279_ (.A(_05300_),
    .B_N(_05301_),
    .X(_05344_));
 sky130_fd_sc_hd__a2bb2o_1 _10280_ (.A1_N(_04901_),
    .A2_N(_05120_),
    .B1(_05298_),
    .B2(_05299_),
    .X(_05345_));
 sky130_fd_sc_hd__a21bo_1 _10281_ (.A1(_04904_),
    .A2(_05221_),
    .B1_N(_05299_),
    .X(_05346_));
 sky130_fd_sc_hd__o21a_1 _10282_ (.A1(_05169_),
    .A2(_05299_),
    .B1(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__xnor2_1 _10283_ (.A(_05345_),
    .B(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__nor2_1 _10284_ (.A(_05344_),
    .B(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__and2_1 _10285_ (.A(_05344_),
    .B(_05348_),
    .X(_05350_));
 sky130_fd_sc_hd__nor2_1 _10286_ (.A(_05349_),
    .B(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__o21a_1 _10287_ (.A1(_05297_),
    .A2(_05225_),
    .B1(_05302_),
    .X(_05352_));
 sky130_fd_sc_hd__a31o_1 _10288_ (.A1(_05227_),
    .A2(_05229_),
    .A3(_05303_),
    .B1(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__xor2_1 _10289_ (.A(_05351_),
    .B(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__xnor2_1 _10290_ (.A(net109),
    .B(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__nor2_1 _10291_ (.A(_05343_),
    .B(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__and2_1 _10292_ (.A(_05343_),
    .B(_05355_),
    .X(_05357_));
 sky130_fd_sc_hd__nor2_1 _10293_ (.A(_05356_),
    .B(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__o21ai_1 _10294_ (.A1(_05341_),
    .A2(_05342_),
    .B1(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__inv_2 _10295_ (.A(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__nor3_1 _10296_ (.A(_05341_),
    .B(_05342_),
    .C(_05358_),
    .Y(_05361_));
 sky130_fd_sc_hd__a211oi_1 _10297_ (.A1(_05340_),
    .A2(_05311_),
    .B1(_05360_),
    .C1(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__o211a_1 _10298_ (.A1(_05360_),
    .A2(_05361_),
    .B1(_05340_),
    .C1(_05311_),
    .X(_05363_));
 sky130_fd_sc_hd__or3_1 _10299_ (.A(_04687_),
    .B(_05362_),
    .C(_05363_),
    .X(_05364_));
 sky130_fd_sc_hd__o21ai_4 _10300_ (.A1(_05337_),
    .A2(_05339_),
    .B1(_05364_),
    .Y(net144));
 sky130_fd_sc_hd__or3_1 _10301_ (.A(_05331_),
    .B(_05332_),
    .C(_05335_),
    .X(_05365_));
 sky130_fd_sc_hd__or2_1 _10302_ (.A(net38),
    .B(net6),
    .X(_05366_));
 sky130_fd_sc_hd__nand2_1 _10303_ (.A(net38),
    .B(net6),
    .Y(_05367_));
 sky130_fd_sc_hd__nand2_1 _10304_ (.A(_05366_),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__xor2_1 _10305_ (.A(_04810_),
    .B(net284),
    .X(_05369_));
 sky130_fd_sc_hd__nor2_1 _10306_ (.A(net92),
    .B(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__inv_2 _10307_ (.A(_04807_),
    .Y(_05371_));
 sky130_fd_sc_hd__o21a_1 _10308_ (.A1(_05371_),
    .A2(net92),
    .B1(_05369_),
    .X(_05372_));
 sky130_fd_sc_hd__a21oi_1 _10309_ (.A1(_04807_),
    .A2(_05370_),
    .B1(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__or3_1 _10310_ (.A(_05320_),
    .B(_05319_),
    .C(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__o21ai_1 _10311_ (.A1(_05320_),
    .A2(_05319_),
    .B1(_05373_),
    .Y(_05375_));
 sky130_fd_sc_hd__nand2_1 _10312_ (.A(_05374_),
    .B(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__a21o_1 _10313_ (.A1(_05323_),
    .A2(_05326_),
    .B1(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__nand3_1 _10314_ (.A(_05323_),
    .B(_05326_),
    .C(_05376_),
    .Y(_05378_));
 sky130_fd_sc_hd__and2_2 _10315_ (.A(_05377_),
    .B(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__xor2_1 _10316_ (.A(_05368_),
    .B(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__a21boi_1 _10317_ (.A1(_05315_),
    .A2(_05328_),
    .B1_N(_05316_),
    .Y(_05381_));
 sky130_fd_sc_hd__xor2_1 _10318_ (.A(_05380_),
    .B(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__nand2_1 _10319_ (.A(_05331_),
    .B(_05382_),
    .Y(_05383_));
 sky130_fd_sc_hd__or2_1 _10320_ (.A(_05331_),
    .B(_05382_),
    .X(_05384_));
 sky130_fd_sc_hd__nand2_1 _10321_ (.A(_05383_),
    .B(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hd__nand3_1 _10322_ (.A(_05365_),
    .B(_05338_),
    .C(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__a21o_1 _10323_ (.A1(_05365_),
    .A2(_05338_),
    .B1(_05385_),
    .X(_05387_));
 sky130_fd_sc_hd__nand2_1 _10324_ (.A(net109),
    .B(_05354_),
    .Y(_05388_));
 sky130_fd_sc_hd__a31o_1 _10325_ (.A1(_05227_),
    .A2(_05229_),
    .A3(_05303_),
    .B1(_05352_),
    .X(_05389_));
 sky130_fd_sc_hd__a21oi_1 _10326_ (.A1(_05351_),
    .A2(_05389_),
    .B1(_05349_),
    .Y(_05390_));
 sky130_fd_sc_hd__nand2_2 _10327_ (.A(_05345_),
    .B(_05347_),
    .Y(_05391_));
 sky130_fd_sc_hd__inv_2 _10328_ (.A(_05222_),
    .Y(_05392_));
 sky130_fd_sc_hd__nor2_1 _10329_ (.A(_05392_),
    .B(_05346_),
    .Y(_05393_));
 sky130_fd_sc_hd__and2_1 _10330_ (.A(_05392_),
    .B(_05346_),
    .X(_05394_));
 sky130_fd_sc_hd__or2_1 _10331_ (.A(_05393_),
    .B(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__xor2_2 _10332_ (.A(_05391_),
    .B(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__xnor2_1 _10333_ (.A(_05390_),
    .B(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__or2_1 _10334_ (.A(net110),
    .B(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__nand2_2 _10335_ (.A(net110),
    .B(_05397_),
    .Y(_05399_));
 sky130_fd_sc_hd__nand2_1 _10336_ (.A(_05398_),
    .B(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__xor2_1 _10337_ (.A(_05388_),
    .B(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__xnor2_1 _10338_ (.A(_05356_),
    .B(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__and2_1 _10339_ (.A(_05340_),
    .B(_05359_),
    .X(_05403_));
 sky130_fd_sc_hd__a21o_1 _10340_ (.A1(_05311_),
    .A2(_05403_),
    .B1(net209),
    .X(_05404_));
 sky130_fd_sc_hd__nand2_1 _10341_ (.A(_05402_),
    .B(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__or2_1 _10342_ (.A(_05402_),
    .B(_05404_),
    .X(_05406_));
 sky130_fd_sc_hd__and3_1 _10343_ (.A(_04463_),
    .B(_05405_),
    .C(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__a31o_4 _10344_ (.A1(_04444_),
    .A2(_05386_),
    .A3(_05387_),
    .B1(_05407_),
    .X(net145));
 sky130_fd_sc_hd__nand2_1 _10345_ (.A(_05356_),
    .B(_05401_),
    .Y(_05408_));
 sky130_fd_sc_hd__or2_1 _10346_ (.A(_05388_),
    .B(_05400_),
    .X(_05409_));
 sky130_fd_sc_hd__o21ai_1 _10347_ (.A1(_05392_),
    .A2(_05346_),
    .B1(_05299_),
    .Y(_05410_));
 sky130_fd_sc_hd__inv_2 _10348_ (.A(_05391_),
    .Y(_05411_));
 sky130_fd_sc_hd__o21ba_1 _10349_ (.A1(_05411_),
    .A2(_05349_),
    .B1_N(_05395_),
    .X(_05412_));
 sky130_fd_sc_hd__a31o_1 _10350_ (.A1(_05351_),
    .A2(_05353_),
    .A3(_05396_),
    .B1(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__xnor2_1 _10351_ (.A(_05410_),
    .B(_05413_),
    .Y(_05414_));
 sky130_fd_sc_hd__or2_1 _10352_ (.A(net111),
    .B(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__nand2_1 _10353_ (.A(net111),
    .B(_05414_),
    .Y(_05416_));
 sky130_fd_sc_hd__nand2_2 _10354_ (.A(_05415_),
    .B(_05416_),
    .Y(_05417_));
 sky130_fd_sc_hd__xor2_2 _10355_ (.A(_05399_),
    .B(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__xor2_2 _10356_ (.A(_05409_),
    .B(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__a21oi_2 _10357_ (.A1(_05408_),
    .A2(_05406_),
    .B1(_05419_),
    .Y(_05420_));
 sky130_fd_sc_hd__a31o_1 _10358_ (.A1(_05408_),
    .A2(_05406_),
    .A3(_05419_),
    .B1(_04688_),
    .X(_05421_));
 sky130_fd_sc_hd__nor2_1 _10359_ (.A(_05380_),
    .B(_05381_),
    .Y(_05422_));
 sky130_fd_sc_hd__or2_1 _10360_ (.A(net39),
    .B(net7),
    .X(_05423_));
 sky130_fd_sc_hd__nand2_1 _10361_ (.A(net39),
    .B(net7),
    .Y(_05424_));
 sky130_fd_sc_hd__nand2_1 _10362_ (.A(_05423_),
    .B(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__xor2_1 _10363_ (.A(net66),
    .B(_04780_),
    .X(_05426_));
 sky130_fd_sc_hd__nor2_1 _10364_ (.A(net284),
    .B(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__inv_2 _10365_ (.A(_04810_),
    .Y(_05428_));
 sky130_fd_sc_hd__o21a_1 _10366_ (.A1(_05428_),
    .A2(net284),
    .B1(_05426_),
    .X(_05429_));
 sky130_fd_sc_hd__a21oi_1 _10367_ (.A1(_04810_),
    .A2(_05427_),
    .B1(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__or3_1 _10368_ (.A(_05371_),
    .B(_05370_),
    .C(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__o21ai_1 _10369_ (.A1(_05371_),
    .A2(_05370_),
    .B1(_05430_),
    .Y(_05432_));
 sky130_fd_sc_hd__nand2_1 _10370_ (.A(_05431_),
    .B(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__a21o_1 _10371_ (.A1(_05374_),
    .A2(_05377_),
    .B1(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__nand3_1 _10372_ (.A(_05374_),
    .B(_05377_),
    .C(_05433_),
    .Y(_05435_));
 sky130_fd_sc_hd__and2_2 _10373_ (.A(_05434_),
    .B(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__xor2_1 _10374_ (.A(_05425_),
    .B(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__a21boi_1 _10375_ (.A1(_05366_),
    .A2(_05379_),
    .B1_N(_05367_),
    .Y(_05438_));
 sky130_fd_sc_hd__xor2_1 _10376_ (.A(_05437_),
    .B(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__nand2_1 _10377_ (.A(_05422_),
    .B(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__or2_1 _10378_ (.A(_05422_),
    .B(_05439_),
    .X(_05441_));
 sky130_fd_sc_hd__nand2_1 _10379_ (.A(_05440_),
    .B(_05441_),
    .Y(_05442_));
 sky130_fd_sc_hd__and3_1 _10380_ (.A(_05383_),
    .B(_05387_),
    .C(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__a21o_1 _10381_ (.A1(_05383_),
    .A2(_05387_),
    .B1(_05442_),
    .X(_05444_));
 sky130_fd_sc_hd__nand2_1 _10382_ (.A(_04724_),
    .B(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__o22ai_4 _10383_ (.A1(_05420_),
    .A2(_05421_),
    .B1(_05443_),
    .B2(_05445_),
    .Y(net146));
 sky130_fd_sc_hd__nor2_1 _10384_ (.A(_05437_),
    .B(_05438_),
    .Y(_05446_));
 sky130_fd_sc_hd__or2_1 _10385_ (.A(net40),
    .B(net8),
    .X(_05447_));
 sky130_fd_sc_hd__nand2_1 _10386_ (.A(net40),
    .B(net8),
    .Y(_05448_));
 sky130_fd_sc_hd__nand2_1 _10387_ (.A(_05447_),
    .B(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__xor2_1 _10388_ (.A(_04814_),
    .B(_04807_),
    .X(_05450_));
 sky130_fd_sc_hd__nor2_1 _10389_ (.A(_04780_),
    .B(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__inv_2 _10390_ (.A(net66),
    .Y(_05452_));
 sky130_fd_sc_hd__o21a_1 _10391_ (.A1(_05452_),
    .A2(_04780_),
    .B1(_05450_),
    .X(_05453_));
 sky130_fd_sc_hd__a21oi_1 _10392_ (.A1(net66),
    .A2(_05451_),
    .B1(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__or3_1 _10393_ (.A(_05428_),
    .B(_05427_),
    .C(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__o21ai_1 _10394_ (.A1(_05428_),
    .A2(_05427_),
    .B1(_05454_),
    .Y(_05456_));
 sky130_fd_sc_hd__nand2_1 _10395_ (.A(_05455_),
    .B(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__a21o_1 _10396_ (.A1(_05431_),
    .A2(_05434_),
    .B1(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__nand3_1 _10397_ (.A(_05431_),
    .B(_05434_),
    .C(_05457_),
    .Y(_05459_));
 sky130_fd_sc_hd__and2_2 _10398_ (.A(_05458_),
    .B(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__xor2_1 _10399_ (.A(_05449_),
    .B(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__a21boi_1 _10400_ (.A1(_05423_),
    .A2(_05436_),
    .B1_N(_05424_),
    .Y(_05462_));
 sky130_fd_sc_hd__xor2_1 _10401_ (.A(_05461_),
    .B(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__nand2_1 _10402_ (.A(_05446_),
    .B(_05463_),
    .Y(_05464_));
 sky130_fd_sc_hd__or2_1 _10403_ (.A(_05446_),
    .B(_05463_),
    .X(_05465_));
 sky130_fd_sc_hd__nand2_1 _10404_ (.A(_05464_),
    .B(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__and3_1 _10405_ (.A(_05440_),
    .B(_05444_),
    .C(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__a21o_1 _10406_ (.A1(_05440_),
    .A2(_05444_),
    .B1(_05466_),
    .X(_05468_));
 sky130_fd_sc_hd__nand2_1 _10407_ (.A(_04724_),
    .B(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__a21bo_1 _10408_ (.A1(_05409_),
    .A2(_05408_),
    .B1_N(_05418_),
    .X(_05470_));
 sky130_fd_sc_hd__a2111o_1 _10409_ (.A1(_05311_),
    .A2(_05403_),
    .B1(_05419_),
    .C1(net209),
    .D1(_05402_),
    .X(_05471_));
 sky130_fd_sc_hd__and2_1 _10410_ (.A(_05470_),
    .B(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__a21o_1 _10411_ (.A1(_05299_),
    .A2(_05413_),
    .B1(_05393_),
    .X(_05473_));
 sky130_fd_sc_hd__xnor2_1 _10412_ (.A(net112),
    .B(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__nand2_1 _10413_ (.A(_05416_),
    .B(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__or2_1 _10414_ (.A(_05416_),
    .B(_05474_),
    .X(_05476_));
 sky130_fd_sc_hd__and2_1 _10415_ (.A(_05475_),
    .B(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__o21bai_1 _10416_ (.A1(_05399_),
    .A2(_05417_),
    .B1_N(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hd__inv_2 _10417_ (.A(net110),
    .Y(_05479_));
 sky130_fd_sc_hd__a21o_1 _10418_ (.A1(_05351_),
    .A2(_05353_),
    .B1(_05349_),
    .X(_05480_));
 sky130_fd_sc_hd__xnor2_1 _10419_ (.A(_05396_),
    .B(_05480_),
    .Y(_05481_));
 sky130_fd_sc_hd__or4b_2 _10420_ (.A(_05479_),
    .B(_05481_),
    .C(_05417_),
    .D_N(_05477_),
    .X(_05482_));
 sky130_fd_sc_hd__nand2_1 _10421_ (.A(_05478_),
    .B(_05482_),
    .Y(_05483_));
 sky130_fd_sc_hd__or2_1 _10422_ (.A(_05472_),
    .B(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__buf_6 _10423_ (.A(_04687_),
    .X(_05485_));
 sky130_fd_sc_hd__a21oi_1 _10424_ (.A1(_05472_),
    .A2(_05483_),
    .B1(_05485_),
    .Y(_05486_));
 sky130_fd_sc_hd__a2bb2o_4 _10425_ (.A1_N(_05467_),
    .A2_N(_05469_),
    .B1(_05484_),
    .B2(_05486_),
    .X(net147));
 sky130_fd_sc_hd__and2_1 _10426_ (.A(net112),
    .B(_05473_),
    .X(_05487_));
 sky130_fd_sc_hd__xnor2_1 _10427_ (.A(net113),
    .B(_05487_),
    .Y(_05488_));
 sky130_fd_sc_hd__xnor2_1 _10428_ (.A(_05476_),
    .B(_05488_),
    .Y(_05489_));
 sky130_fd_sc_hd__a21oi_1 _10429_ (.A1(_05482_),
    .A2(_05484_),
    .B1(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__a31o_1 _10430_ (.A1(_05482_),
    .A2(_05484_),
    .A3(_05489_),
    .B1(_04688_),
    .X(_05491_));
 sky130_fd_sc_hd__nor2_1 _10431_ (.A(_05461_),
    .B(_05462_),
    .Y(_05492_));
 sky130_fd_sc_hd__or2_1 _10432_ (.A(net41),
    .B(net9),
    .X(_05493_));
 sky130_fd_sc_hd__nand2_1 _10433_ (.A(net41),
    .B(net9),
    .Y(_05494_));
 sky130_fd_sc_hd__nand2_1 _10434_ (.A(_05493_),
    .B(_05494_),
    .Y(_05495_));
 sky130_fd_sc_hd__xor2_1 _10435_ (.A(net68),
    .B(_04810_),
    .X(_05496_));
 sky130_fd_sc_hd__nor2_1 _10436_ (.A(_04807_),
    .B(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__inv_2 _10437_ (.A(_04814_),
    .Y(_05498_));
 sky130_fd_sc_hd__o21a_1 _10438_ (.A1(_05498_),
    .A2(_04807_),
    .B1(_05496_),
    .X(_05499_));
 sky130_fd_sc_hd__a21oi_1 _10439_ (.A1(_04814_),
    .A2(_05497_),
    .B1(_05499_),
    .Y(_05500_));
 sky130_fd_sc_hd__or3_1 _10440_ (.A(_05452_),
    .B(_05451_),
    .C(_05500_),
    .X(_05501_));
 sky130_fd_sc_hd__o21ai_1 _10441_ (.A1(_05452_),
    .A2(_05451_),
    .B1(_05500_),
    .Y(_05502_));
 sky130_fd_sc_hd__nand2_1 _10442_ (.A(_05501_),
    .B(_05502_),
    .Y(_05503_));
 sky130_fd_sc_hd__a21o_1 _10443_ (.A1(_05455_),
    .A2(_05458_),
    .B1(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__nand3_1 _10444_ (.A(_05455_),
    .B(_05458_),
    .C(_05503_),
    .Y(_05505_));
 sky130_fd_sc_hd__and2_2 _10445_ (.A(_05504_),
    .B(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__xor2_1 _10446_ (.A(_05495_),
    .B(_05506_),
    .X(_05507_));
 sky130_fd_sc_hd__a21boi_1 _10447_ (.A1(_05447_),
    .A2(_05460_),
    .B1_N(_05448_),
    .Y(_05508_));
 sky130_fd_sc_hd__xor2_1 _10448_ (.A(_05507_),
    .B(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__nand2_1 _10449_ (.A(_05492_),
    .B(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__or2_1 _10450_ (.A(_05492_),
    .B(_05509_),
    .X(_05511_));
 sky130_fd_sc_hd__nand2_1 _10451_ (.A(_05510_),
    .B(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__and3_1 _10452_ (.A(_05464_),
    .B(_05468_),
    .C(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__a21o_1 _10453_ (.A1(_05464_),
    .A2(_05468_),
    .B1(_05512_),
    .X(_05514_));
 sky130_fd_sc_hd__nand2_1 _10454_ (.A(_04724_),
    .B(_05514_),
    .Y(_05515_));
 sky130_fd_sc_hd__o22ai_1 _10455_ (.A1(_05490_),
    .A2(_05491_),
    .B1(_05513_),
    .B2(_05515_),
    .Y(net148));
 sky130_fd_sc_hd__nor2_1 _10456_ (.A(_05507_),
    .B(_05508_),
    .Y(_05516_));
 sky130_fd_sc_hd__or2_1 _10457_ (.A(net42),
    .B(net10),
    .X(_05517_));
 sky130_fd_sc_hd__nand2_1 _10458_ (.A(net42),
    .B(net10),
    .Y(_05518_));
 sky130_fd_sc_hd__nand2_1 _10459_ (.A(_05517_),
    .B(_05518_),
    .Y(_05519_));
 sky130_fd_sc_hd__xor2_1 _10460_ (.A(net69),
    .B(net66),
    .X(_05520_));
 sky130_fd_sc_hd__nor2_1 _10461_ (.A(_04810_),
    .B(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__inv_2 _10462_ (.A(net68),
    .Y(_05522_));
 sky130_fd_sc_hd__o21a_1 _10463_ (.A1(_05522_),
    .A2(_04810_),
    .B1(_05520_),
    .X(_05523_));
 sky130_fd_sc_hd__a21oi_1 _10464_ (.A1(net68),
    .A2(_05521_),
    .B1(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__or3_1 _10465_ (.A(_05498_),
    .B(_05497_),
    .C(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__o21ai_1 _10466_ (.A1(_05498_),
    .A2(_05497_),
    .B1(_05524_),
    .Y(_05526_));
 sky130_fd_sc_hd__nand2_1 _10467_ (.A(_05525_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__a21o_1 _10468_ (.A1(_05501_),
    .A2(_05504_),
    .B1(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__nand3_1 _10469_ (.A(_05501_),
    .B(_05504_),
    .C(_05527_),
    .Y(_05529_));
 sky130_fd_sc_hd__and2_2 _10470_ (.A(_05528_),
    .B(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__xor2_1 _10471_ (.A(_05519_),
    .B(_05530_),
    .X(_05531_));
 sky130_fd_sc_hd__a21boi_1 _10472_ (.A1(_05493_),
    .A2(_05506_),
    .B1_N(_05494_),
    .Y(_05532_));
 sky130_fd_sc_hd__xor2_1 _10473_ (.A(_05531_),
    .B(_05532_),
    .X(_05533_));
 sky130_fd_sc_hd__nand2_1 _10474_ (.A(_05516_),
    .B(_05533_),
    .Y(_05534_));
 sky130_fd_sc_hd__or2_1 _10475_ (.A(_05516_),
    .B(_05533_),
    .X(_05535_));
 sky130_fd_sc_hd__nand2_1 _10476_ (.A(_05534_),
    .B(_05535_),
    .Y(_05536_));
 sky130_fd_sc_hd__and3_1 _10477_ (.A(_05510_),
    .B(_05514_),
    .C(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__a21o_1 _10478_ (.A1(_05510_),
    .A2(_05514_),
    .B1(_05536_),
    .X(_05538_));
 sky130_fd_sc_hd__nand2_1 _10479_ (.A(_04724_),
    .B(_05538_),
    .Y(_05539_));
 sky130_fd_sc_hd__and3_1 _10480_ (.A(net113),
    .B(net114),
    .C(_05487_),
    .X(_05540_));
 sky130_fd_sc_hd__a31o_1 _10481_ (.A1(net112),
    .A2(net113),
    .A3(_05473_),
    .B1(net114),
    .X(_05541_));
 sky130_fd_sc_hd__or2b_1 _10482_ (.A(_05540_),
    .B_N(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__a211o_1 _10483_ (.A1(_05470_),
    .A2(_05471_),
    .B1(_05483_),
    .C1(_05489_),
    .X(_05543_));
 sky130_fd_sc_hd__a21o_1 _10484_ (.A1(_05476_),
    .A2(_05482_),
    .B1(_05488_),
    .X(_05544_));
 sky130_fd_sc_hd__and3_1 _10485_ (.A(_05542_),
    .B(_05543_),
    .C(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__a21oi_2 _10486_ (.A1(_05543_),
    .A2(_05544_),
    .B1(_05542_),
    .Y(_05546_));
 sky130_fd_sc_hd__or3_1 _10487_ (.A(_04687_),
    .B(_05545_),
    .C(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__o21ai_4 _10488_ (.A1(_05537_),
    .A2(_05539_),
    .B1(_05547_),
    .Y(net149));
 sky130_fd_sc_hd__nor2_1 _10489_ (.A(_05531_),
    .B(_05532_),
    .Y(_05548_));
 sky130_fd_sc_hd__or2_1 _10490_ (.A(net43),
    .B(net11),
    .X(_05549_));
 sky130_fd_sc_hd__nand2_1 _10491_ (.A(net43),
    .B(net11),
    .Y(_05550_));
 sky130_fd_sc_hd__nand2_1 _10492_ (.A(_05549_),
    .B(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__xor2_1 _10493_ (.A(net70),
    .B(_04814_),
    .X(_05552_));
 sky130_fd_sc_hd__nor2_1 _10494_ (.A(net66),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__inv_2 _10495_ (.A(net69),
    .Y(_05554_));
 sky130_fd_sc_hd__o21a_1 _10496_ (.A1(_05554_),
    .A2(net66),
    .B1(_05552_),
    .X(_05555_));
 sky130_fd_sc_hd__a21oi_2 _10497_ (.A1(net69),
    .A2(_05553_),
    .B1(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__or3_2 _10498_ (.A(_05522_),
    .B(_05521_),
    .C(_05556_),
    .X(_05557_));
 sky130_fd_sc_hd__o21ai_1 _10499_ (.A1(_05522_),
    .A2(_05521_),
    .B1(_05556_),
    .Y(_05558_));
 sky130_fd_sc_hd__nand2_1 _10500_ (.A(_05557_),
    .B(_05558_),
    .Y(_05559_));
 sky130_fd_sc_hd__a21o_1 _10501_ (.A1(_05525_),
    .A2(_05528_),
    .B1(_05559_),
    .X(_05560_));
 sky130_fd_sc_hd__nand3_1 _10502_ (.A(_05525_),
    .B(_05528_),
    .C(_05559_),
    .Y(_05561_));
 sky130_fd_sc_hd__and2_2 _10503_ (.A(_05560_),
    .B(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__xor2_1 _10504_ (.A(_05551_),
    .B(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__a21boi_1 _10505_ (.A1(_05517_),
    .A2(_05530_),
    .B1_N(_05518_),
    .Y(_05564_));
 sky130_fd_sc_hd__xor2_1 _10506_ (.A(_05563_),
    .B(_05564_),
    .X(_05565_));
 sky130_fd_sc_hd__nand2_1 _10507_ (.A(_05548_),
    .B(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__or2_1 _10508_ (.A(_05548_),
    .B(_05565_),
    .X(_05567_));
 sky130_fd_sc_hd__nand2_1 _10509_ (.A(_05566_),
    .B(_05567_),
    .Y(_05568_));
 sky130_fd_sc_hd__and3_1 _10510_ (.A(_05534_),
    .B(_05538_),
    .C(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__a21o_1 _10511_ (.A1(_05534_),
    .A2(_05538_),
    .B1(_05568_),
    .X(_05570_));
 sky130_fd_sc_hd__nand2_1 _10512_ (.A(_04724_),
    .B(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__or2_1 _10513_ (.A(_05540_),
    .B(_05546_),
    .X(_05572_));
 sky130_fd_sc_hd__nand2_1 _10514_ (.A(net115),
    .B(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__o21a_1 _10515_ (.A1(net115),
    .A2(_05572_),
    .B1(_04463_),
    .X(_05574_));
 sky130_fd_sc_hd__a2bb2o_4 _10516_ (.A1_N(_05569_),
    .A2_N(_05571_),
    .B1(_05573_),
    .B2(_05574_),
    .X(net150));
 sky130_fd_sc_hd__nor2_1 _10517_ (.A(_05563_),
    .B(_05564_),
    .Y(_05575_));
 sky130_fd_sc_hd__or2_1 _10518_ (.A(net45),
    .B(net13),
    .X(_05576_));
 sky130_fd_sc_hd__nand2_1 _10519_ (.A(net45),
    .B(net13),
    .Y(_05577_));
 sky130_fd_sc_hd__nand2_1 _10520_ (.A(_05576_),
    .B(_05577_),
    .Y(_05578_));
 sky130_fd_sc_hd__xor2_1 _10521_ (.A(_04826_),
    .B(net68),
    .X(_05579_));
 sky130_fd_sc_hd__nor2_1 _10522_ (.A(_04814_),
    .B(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__o21a_1 _10523_ (.A1(_04828_),
    .A2(_04814_),
    .B1(_05579_),
    .X(_05581_));
 sky130_fd_sc_hd__a21oi_1 _10524_ (.A1(net70),
    .A2(_05580_),
    .B1(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__or3_1 _10525_ (.A(_05554_),
    .B(_05553_),
    .C(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__o21ai_1 _10526_ (.A1(_05554_),
    .A2(_05553_),
    .B1(_05582_),
    .Y(_05584_));
 sky130_fd_sc_hd__nand2_1 _10527_ (.A(_05583_),
    .B(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__a21o_1 _10528_ (.A1(_05557_),
    .A2(_05560_),
    .B1(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__nand3_1 _10529_ (.A(_05557_),
    .B(_05560_),
    .C(_05585_),
    .Y(_05587_));
 sky130_fd_sc_hd__and2_2 _10530_ (.A(_05586_),
    .B(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__xor2_1 _10531_ (.A(_05578_),
    .B(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__a21boi_1 _10532_ (.A1(_05549_),
    .A2(_05562_),
    .B1_N(_05550_),
    .Y(_05590_));
 sky130_fd_sc_hd__xor2_1 _10533_ (.A(_05589_),
    .B(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__nand2_1 _10534_ (.A(_05575_),
    .B(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__or2_1 _10535_ (.A(_05575_),
    .B(_05591_),
    .X(_05593_));
 sky130_fd_sc_hd__nand2_1 _10536_ (.A(_05592_),
    .B(_05593_),
    .Y(_05594_));
 sky130_fd_sc_hd__and3_1 _10537_ (.A(_05566_),
    .B(_05570_),
    .C(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__a21o_1 _10538_ (.A1(_05566_),
    .A2(_05570_),
    .B1(_05594_),
    .X(_05596_));
 sky130_fd_sc_hd__nand2_1 _10539_ (.A(_04724_),
    .B(_05596_),
    .Y(_05597_));
 sky130_fd_sc_hd__inv_2 _10540_ (.A(net117),
    .Y(_05598_));
 sky130_fd_sc_hd__nor2_1 _10541_ (.A(_05598_),
    .B(_05573_),
    .Y(_05599_));
 sky130_fd_sc_hd__a21o_1 _10542_ (.A1(_05598_),
    .A2(_05573_),
    .B1(_04688_),
    .X(_05600_));
 sky130_fd_sc_hd__o22ai_4 _10543_ (.A1(_05595_),
    .A2(_05597_),
    .B1(_05599_),
    .B2(_05600_),
    .Y(net152));
 sky130_fd_sc_hd__nor2_1 _10544_ (.A(_05589_),
    .B(_05590_),
    .Y(_05601_));
 sky130_fd_sc_hd__xor2_1 _10545_ (.A(net72),
    .B(net69),
    .X(_05602_));
 sky130_fd_sc_hd__nor2_1 _10546_ (.A(net68),
    .B(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__inv_2 _10547_ (.A(_04826_),
    .Y(_05604_));
 sky130_fd_sc_hd__o21a_1 _10548_ (.A1(_05604_),
    .A2(net68),
    .B1(_05602_),
    .X(_05605_));
 sky130_fd_sc_hd__a21oi_1 _10549_ (.A1(_04826_),
    .A2(_05603_),
    .B1(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__or3_1 _10550_ (.A(_04828_),
    .B(_05580_),
    .C(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__o21ai_1 _10551_ (.A1(_04828_),
    .A2(_05580_),
    .B1(_05606_),
    .Y(_05608_));
 sky130_fd_sc_hd__nand2_1 _10552_ (.A(_05607_),
    .B(_05608_),
    .Y(_05609_));
 sky130_fd_sc_hd__a21o_1 _10553_ (.A1(_05583_),
    .A2(_05586_),
    .B1(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__nand3_1 _10554_ (.A(_05583_),
    .B(_05586_),
    .C(_05609_),
    .Y(_05611_));
 sky130_fd_sc_hd__and2_1 _10555_ (.A(_05610_),
    .B(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__nor2_1 _10556_ (.A(net46),
    .B(net14),
    .Y(_05613_));
 sky130_fd_sc_hd__and2_1 _10557_ (.A(net46),
    .B(net14),
    .X(_05614_));
 sky130_fd_sc_hd__nor2_1 _10558_ (.A(_05613_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__xnor2_1 _10559_ (.A(_05612_),
    .B(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__a21bo_1 _10560_ (.A1(_05576_),
    .A2(_05588_),
    .B1_N(_05577_),
    .X(_05617_));
 sky130_fd_sc_hd__xnor2_1 _10561_ (.A(_05616_),
    .B(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand2_1 _10562_ (.A(_05601_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__or2_1 _10563_ (.A(_05601_),
    .B(_05618_),
    .X(_05620_));
 sky130_fd_sc_hd__nand2_1 _10564_ (.A(_05619_),
    .B(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__and3_1 _10565_ (.A(_05592_),
    .B(_05596_),
    .C(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__a21o_1 _10566_ (.A1(_05592_),
    .A2(_05596_),
    .B1(_05621_),
    .X(_05623_));
 sky130_fd_sc_hd__nand2_1 _10567_ (.A(_04724_),
    .B(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__o2111ai_4 _10568_ (.A1(_05540_),
    .A2(_05546_),
    .B1(net115),
    .C1(net117),
    .D1(net118),
    .Y(_05625_));
 sky130_fd_sc_hd__o21a_1 _10569_ (.A1(net118),
    .A2(_05599_),
    .B1(_04463_),
    .X(_05626_));
 sky130_fd_sc_hd__a2bb2o_4 _10570_ (.A1_N(_05622_),
    .A2_N(_05624_),
    .B1(_05625_),
    .B2(_05626_),
    .X(net153));
 sky130_fd_sc_hd__nand2_1 _10571_ (.A(_05619_),
    .B(_05623_),
    .Y(_05627_));
 sky130_fd_sc_hd__or2b_1 _10572_ (.A(_05616_),
    .B_N(_05617_),
    .X(_05628_));
 sky130_fd_sc_hd__or2_1 _10573_ (.A(net47),
    .B(net15),
    .X(_05629_));
 sky130_fd_sc_hd__nand2_1 _10574_ (.A(net47),
    .B(net15),
    .Y(_05630_));
 sky130_fd_sc_hd__nand2_1 _10575_ (.A(_05629_),
    .B(_05630_),
    .Y(_05631_));
 sky130_fd_sc_hd__xor2_1 _10576_ (.A(_04770_),
    .B(net70),
    .X(_05632_));
 sky130_fd_sc_hd__nor2_1 _10577_ (.A(net69),
    .B(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__o21a_1 _10578_ (.A1(_04766_),
    .A2(net69),
    .B1(_05632_),
    .X(_05634_));
 sky130_fd_sc_hd__a21oi_1 _10579_ (.A1(net72),
    .A2(_05633_),
    .B1(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__or3_1 _10580_ (.A(_05604_),
    .B(_05603_),
    .C(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__o21ai_1 _10581_ (.A1(_05604_),
    .A2(_05603_),
    .B1(_05635_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand2_1 _10582_ (.A(_05636_),
    .B(_05637_),
    .Y(_05638_));
 sky130_fd_sc_hd__a21o_1 _10583_ (.A1(_05607_),
    .A2(_05610_),
    .B1(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__nand3_1 _10584_ (.A(_05607_),
    .B(_05610_),
    .C(_05638_),
    .Y(_05640_));
 sky130_fd_sc_hd__and2_1 _10585_ (.A(_05639_),
    .B(_05640_),
    .X(_05641_));
 sky130_fd_sc_hd__xor2_1 _10586_ (.A(_05631_),
    .B(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__a21oi_1 _10587_ (.A1(_05612_),
    .A2(_05615_),
    .B1(_05614_),
    .Y(_05643_));
 sky130_fd_sc_hd__nor2_1 _10588_ (.A(_05642_),
    .B(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__and2_1 _10589_ (.A(_05642_),
    .B(_05643_),
    .X(_05645_));
 sky130_fd_sc_hd__or2_1 _10590_ (.A(_05644_),
    .B(_05645_),
    .X(_05646_));
 sky130_fd_sc_hd__or2_1 _10591_ (.A(_05628_),
    .B(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__nand2_1 _10592_ (.A(_05628_),
    .B(_05646_),
    .Y(_05648_));
 sky130_fd_sc_hd__nand2_1 _10593_ (.A(_05647_),
    .B(_05648_),
    .Y(_05649_));
 sky130_fd_sc_hd__xor2_1 _10594_ (.A(_05627_),
    .B(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__inv_2 _10595_ (.A(net119),
    .Y(_05651_));
 sky130_fd_sc_hd__or2_1 _10596_ (.A(_05651_),
    .B(_05625_),
    .X(_05652_));
 sky130_fd_sc_hd__a21oi_1 _10597_ (.A1(_05651_),
    .A2(_05625_),
    .B1(_05485_),
    .Y(_05653_));
 sky130_fd_sc_hd__a2bb2o_2 _10598_ (.A1_N(_04956_),
    .A2_N(_05650_),
    .B1(_05652_),
    .B2(_05653_),
    .X(net154));
 sky130_fd_sc_hd__a21bo_1 _10599_ (.A1(_05619_),
    .A2(_05623_),
    .B1_N(_05648_),
    .X(_05654_));
 sky130_fd_sc_hd__or2_1 _10600_ (.A(net48),
    .B(net16),
    .X(_05655_));
 sky130_fd_sc_hd__nand2_1 _10601_ (.A(net48),
    .B(net16),
    .Y(_05656_));
 sky130_fd_sc_hd__nand2_1 _10602_ (.A(_05655_),
    .B(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__xor2_1 _10603_ (.A(net74),
    .B(_04826_),
    .X(_05658_));
 sky130_fd_sc_hd__nor2_1 _10604_ (.A(net70),
    .B(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__inv_2 _10605_ (.A(_04770_),
    .Y(_05660_));
 sky130_fd_sc_hd__o21a_1 _10606_ (.A1(_05660_),
    .A2(net70),
    .B1(_05658_),
    .X(_05661_));
 sky130_fd_sc_hd__a21oi_1 _10607_ (.A1(_04770_),
    .A2(_05659_),
    .B1(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__or3_1 _10608_ (.A(_04766_),
    .B(_05633_),
    .C(_05662_),
    .X(_05663_));
 sky130_fd_sc_hd__o21ai_1 _10609_ (.A1(_04766_),
    .A2(_05633_),
    .B1(_05662_),
    .Y(_05664_));
 sky130_fd_sc_hd__nand2_1 _10610_ (.A(_05663_),
    .B(_05664_),
    .Y(_05665_));
 sky130_fd_sc_hd__a21o_1 _10611_ (.A1(_05636_),
    .A2(_05639_),
    .B1(_05665_),
    .X(_05666_));
 sky130_fd_sc_hd__nand3_1 _10612_ (.A(_05636_),
    .B(_05639_),
    .C(_05665_),
    .Y(_05667_));
 sky130_fd_sc_hd__and2_1 _10613_ (.A(_05666_),
    .B(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__xor2_1 _10614_ (.A(_05657_),
    .B(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__a21boi_1 _10615_ (.A1(_05629_),
    .A2(_05641_),
    .B1_N(_05630_),
    .Y(_05670_));
 sky130_fd_sc_hd__nor2_1 _10616_ (.A(_05669_),
    .B(_05670_),
    .Y(_05671_));
 sky130_fd_sc_hd__and2_1 _10617_ (.A(_05669_),
    .B(_05670_),
    .X(_05672_));
 sky130_fd_sc_hd__nor2_1 _10618_ (.A(_05671_),
    .B(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__or2_1 _10619_ (.A(_05644_),
    .B(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__nand2_1 _10620_ (.A(_05644_),
    .B(_05673_),
    .Y(_05675_));
 sky130_fd_sc_hd__nand2_1 _10621_ (.A(_05674_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__a21oi_1 _10622_ (.A1(_05647_),
    .A2(_05654_),
    .B1(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hd__a31o_1 _10623_ (.A1(_05647_),
    .A2(_05654_),
    .A3(_05676_),
    .B1(_04956_),
    .X(_05678_));
 sky130_fd_sc_hd__xnor2_1 _10624_ (.A(net120),
    .B(_05652_),
    .Y(_05679_));
 sky130_fd_sc_hd__a2bb2o_4 _10625_ (.A1_N(_05677_),
    .A2_N(_05678_),
    .B1(_05679_),
    .B2(_04464_),
    .X(net155));
 sky130_fd_sc_hd__or2_1 _10626_ (.A(net49),
    .B(net17),
    .X(_05680_));
 sky130_fd_sc_hd__nand2_1 _10627_ (.A(net49),
    .B(net17),
    .Y(_05681_));
 sky130_fd_sc_hd__nand2_1 _10628_ (.A(_05680_),
    .B(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__xor2_1 _10629_ (.A(_04773_),
    .B(net72),
    .X(_05683_));
 sky130_fd_sc_hd__nor2_1 _10630_ (.A(_04826_),
    .B(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__o21a_1 _10631_ (.A1(_04775_),
    .A2(_04826_),
    .B1(_05683_),
    .X(_05685_));
 sky130_fd_sc_hd__a21oi_1 _10632_ (.A1(net74),
    .A2(_05684_),
    .B1(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__or3_1 _10633_ (.A(_05660_),
    .B(_05659_),
    .C(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__o21ai_1 _10634_ (.A1(_05660_),
    .A2(_05659_),
    .B1(_05686_),
    .Y(_05688_));
 sky130_fd_sc_hd__nand2_1 _10635_ (.A(_05687_),
    .B(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__a21o_1 _10636_ (.A1(_05663_),
    .A2(_05666_),
    .B1(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__nand3_1 _10637_ (.A(_05663_),
    .B(_05666_),
    .C(_05689_),
    .Y(_05691_));
 sky130_fd_sc_hd__and2_1 _10638_ (.A(_05690_),
    .B(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__xor2_1 _10639_ (.A(_05682_),
    .B(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__a21boi_1 _10640_ (.A1(_05655_),
    .A2(_05668_),
    .B1_N(_05656_),
    .Y(_05694_));
 sky130_fd_sc_hd__xor2_1 _10641_ (.A(_05693_),
    .B(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__nand2_1 _10642_ (.A(_05671_),
    .B(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__or2_1 _10643_ (.A(_05671_),
    .B(_05695_),
    .X(_05697_));
 sky130_fd_sc_hd__nand2_1 _10644_ (.A(_05696_),
    .B(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__a21bo_1 _10645_ (.A1(_05647_),
    .A2(_05654_),
    .B1_N(_05674_),
    .X(_05699_));
 sky130_fd_sc_hd__nand3_1 _10646_ (.A(_05675_),
    .B(_05698_),
    .C(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__a21o_1 _10647_ (.A1(_05675_),
    .A2(_05699_),
    .B1(_05698_),
    .X(_05701_));
 sky130_fd_sc_hd__inv_2 _10648_ (.A(net120),
    .Y(_05702_));
 sky130_fd_sc_hd__inv_2 _10649_ (.A(net121),
    .Y(_05703_));
 sky130_fd_sc_hd__o21a_1 _10650_ (.A1(_05702_),
    .A2(_05652_),
    .B1(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__nor4_1 _10651_ (.A(_05651_),
    .B(_05702_),
    .C(_05703_),
    .D(_05625_),
    .Y(_05705_));
 sky130_fd_sc_hd__nor3_1 _10652_ (.A(_04688_),
    .B(_05704_),
    .C(_05705_),
    .Y(_05706_));
 sky130_fd_sc_hd__a31o_4 _10653_ (.A1(_04444_),
    .A2(_05700_),
    .A3(_05701_),
    .B1(_05706_),
    .X(net156));
 sky130_fd_sc_hd__nor2_1 _10654_ (.A(_05693_),
    .B(_05694_),
    .Y(_05707_));
 sky130_fd_sc_hd__xor2_1 _10655_ (.A(net77),
    .B(_04770_),
    .X(_05708_));
 sky130_fd_sc_hd__nor2_1 _10656_ (.A(net72),
    .B(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__inv_2 _10657_ (.A(_04773_),
    .Y(_05710_));
 sky130_fd_sc_hd__o21a_1 _10658_ (.A1(_05710_),
    .A2(net72),
    .B1(_05708_),
    .X(_05711_));
 sky130_fd_sc_hd__a21oi_1 _10659_ (.A1(_04773_),
    .A2(_05709_),
    .B1(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__or3_1 _10660_ (.A(_04775_),
    .B(_05684_),
    .C(_05712_),
    .X(_05713_));
 sky130_fd_sc_hd__o21ai_1 _10661_ (.A1(_04775_),
    .A2(_05684_),
    .B1(_05712_),
    .Y(_05714_));
 sky130_fd_sc_hd__nand2_1 _10662_ (.A(_05713_),
    .B(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hd__a21o_1 _10663_ (.A1(_05687_),
    .A2(_05690_),
    .B1(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__nand3_1 _10664_ (.A(_05687_),
    .B(_05690_),
    .C(_05715_),
    .Y(_05717_));
 sky130_fd_sc_hd__and2_1 _10665_ (.A(_05716_),
    .B(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__nor2_1 _10666_ (.A(net50),
    .B(net18),
    .Y(_05719_));
 sky130_fd_sc_hd__and2_1 _10667_ (.A(net50),
    .B(net18),
    .X(_05720_));
 sky130_fd_sc_hd__nor2_1 _10668_ (.A(_05719_),
    .B(_05720_),
    .Y(_05721_));
 sky130_fd_sc_hd__xnor2_1 _10669_ (.A(_05718_),
    .B(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__a21bo_1 _10670_ (.A1(_05680_),
    .A2(_05692_),
    .B1_N(_05681_),
    .X(_05723_));
 sky130_fd_sc_hd__xnor2_1 _10671_ (.A(_05722_),
    .B(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__nand2_1 _10672_ (.A(_05707_),
    .B(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__or2_1 _10673_ (.A(_05707_),
    .B(_05724_),
    .X(_05726_));
 sky130_fd_sc_hd__nand2_1 _10674_ (.A(_05725_),
    .B(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__and3_1 _10675_ (.A(_05696_),
    .B(_05701_),
    .C(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__a21o_1 _10676_ (.A1(_05696_),
    .A2(_05701_),
    .B1(_05727_),
    .X(_05729_));
 sky130_fd_sc_hd__nand2_1 _10677_ (.A(_04443_),
    .B(_05729_),
    .Y(_05730_));
 sky130_fd_sc_hd__and2_2 _10678_ (.A(net122),
    .B(net202),
    .X(_05731_));
 sky130_fd_sc_hd__o21ai_1 _10679_ (.A1(net122),
    .A2(net203),
    .B1(_04463_),
    .Y(_05732_));
 sky130_fd_sc_hd__o22ai_4 _10680_ (.A1(_05728_),
    .A2(_05730_),
    .B1(_05731_),
    .B2(_05732_),
    .Y(net157));
 sky130_fd_sc_hd__and2b_1 _10681_ (.A_N(_05722_),
    .B(_05723_),
    .X(_05733_));
 sky130_fd_sc_hd__or2_1 _10682_ (.A(net51),
    .B(net19),
    .X(_05734_));
 sky130_fd_sc_hd__nand2_1 _10683_ (.A(net51),
    .B(net19),
    .Y(_05735_));
 sky130_fd_sc_hd__nand2_1 _10684_ (.A(_05734_),
    .B(_05735_),
    .Y(_05736_));
 sky130_fd_sc_hd__nand2_1 _10685_ (.A(net78),
    .B(_04775_),
    .Y(_05737_));
 sky130_fd_sc_hd__inv_2 _10686_ (.A(net78),
    .Y(_05738_));
 sky130_fd_sc_hd__nand2_1 _10687_ (.A(_05738_),
    .B(net74),
    .Y(_05739_));
 sky130_fd_sc_hd__nand2_1 _10688_ (.A(_05737_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__nor2_1 _10689_ (.A(_04770_),
    .B(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__o21a_1 _10690_ (.A1(_04753_),
    .A2(_04770_),
    .B1(_05740_),
    .X(_05742_));
 sky130_fd_sc_hd__a21oi_1 _10691_ (.A1(net77),
    .A2(_05741_),
    .B1(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__or3_1 _10692_ (.A(_05710_),
    .B(_05709_),
    .C(_05743_),
    .X(_05744_));
 sky130_fd_sc_hd__o21ai_1 _10693_ (.A1(_05710_),
    .A2(_05709_),
    .B1(_05743_),
    .Y(_05745_));
 sky130_fd_sc_hd__nand2_1 _10694_ (.A(_05744_),
    .B(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__a21o_1 _10695_ (.A1(_05713_),
    .A2(_05716_),
    .B1(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__nand3_1 _10696_ (.A(_05713_),
    .B(_05716_),
    .C(_05746_),
    .Y(_05748_));
 sky130_fd_sc_hd__and2_1 _10697_ (.A(_05747_),
    .B(_05748_),
    .X(_05749_));
 sky130_fd_sc_hd__xor2_1 _10698_ (.A(_05736_),
    .B(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__a21oi_1 _10699_ (.A1(_05718_),
    .A2(_05721_),
    .B1(_05720_),
    .Y(_05751_));
 sky130_fd_sc_hd__nor2_1 _10700_ (.A(_05750_),
    .B(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__and2_1 _10701_ (.A(_05750_),
    .B(_05751_),
    .X(_05753_));
 sky130_fd_sc_hd__nor2_1 _10702_ (.A(_05752_),
    .B(_05753_),
    .Y(_05754_));
 sky130_fd_sc_hd__xnor2_1 _10703_ (.A(_05733_),
    .B(_05754_),
    .Y(_05755_));
 sky130_fd_sc_hd__a21oi_1 _10704_ (.A1(_05725_),
    .A2(_05729_),
    .B1(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__a31o_1 _10705_ (.A1(_05725_),
    .A2(_05729_),
    .A3(_05755_),
    .B1(_04956_),
    .X(_05757_));
 sky130_fd_sc_hd__xor2_1 _10706_ (.A(net123),
    .B(_05731_),
    .X(_05758_));
 sky130_fd_sc_hd__a2bb2o_4 _10707_ (.A1_N(_05756_),
    .A2_N(_05757_),
    .B1(_05758_),
    .B2(_04464_),
    .X(net158));
 sky130_fd_sc_hd__a21oi_1 _10708_ (.A1(net123),
    .A2(_05731_),
    .B1(net124),
    .Y(_05759_));
 sky130_fd_sc_hd__and4_2 _10709_ (.A(net122),
    .B(net123),
    .C(net124),
    .D(net202),
    .X(_05760_));
 sky130_fd_sc_hd__nand2_1 _10710_ (.A(_05733_),
    .B(_05754_),
    .Y(_05761_));
 sky130_fd_sc_hd__a21o_1 _10711_ (.A1(_05725_),
    .A2(_05729_),
    .B1(_05755_),
    .X(_05762_));
 sky130_fd_sc_hd__or2_1 _10712_ (.A(net52),
    .B(net20),
    .X(_05763_));
 sky130_fd_sc_hd__nand2_1 _10713_ (.A(net52),
    .B(net20),
    .Y(_05764_));
 sky130_fd_sc_hd__nand2_1 _10714_ (.A(_05763_),
    .B(_05764_),
    .Y(_05765_));
 sky130_fd_sc_hd__or2_1 _10715_ (.A(_04753_),
    .B(_05741_),
    .X(_05766_));
 sky130_fd_sc_hd__xor2_1 _10716_ (.A(net79),
    .B(_04773_),
    .X(_05767_));
 sky130_fd_sc_hd__or2_1 _10717_ (.A(net74),
    .B(_05767_),
    .X(_05768_));
 sky130_fd_sc_hd__o2bb2a_1 _10718_ (.A1_N(_05737_),
    .A2_N(_05767_),
    .B1(_05768_),
    .B2(_05738_),
    .X(_05769_));
 sky130_fd_sc_hd__or2_1 _10719_ (.A(_05766_),
    .B(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__nand2_1 _10720_ (.A(_05766_),
    .B(_05769_),
    .Y(_05771_));
 sky130_fd_sc_hd__nand2_1 _10721_ (.A(_05770_),
    .B(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__a21o_1 _10722_ (.A1(_05744_),
    .A2(_05747_),
    .B1(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__nand3_1 _10723_ (.A(_05744_),
    .B(_05747_),
    .C(_05772_),
    .Y(_05774_));
 sky130_fd_sc_hd__and2_1 _10724_ (.A(_05773_),
    .B(_05774_),
    .X(_05775_));
 sky130_fd_sc_hd__xor2_1 _10725_ (.A(_05765_),
    .B(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__a21boi_1 _10726_ (.A1(_05734_),
    .A2(_05749_),
    .B1_N(_05735_),
    .Y(_05777_));
 sky130_fd_sc_hd__nor2_1 _10727_ (.A(_05776_),
    .B(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__and2_1 _10728_ (.A(_05776_),
    .B(_05777_),
    .X(_05779_));
 sky130_fd_sc_hd__nor2_1 _10729_ (.A(_05778_),
    .B(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__xnor2_1 _10730_ (.A(_05752_),
    .B(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__a21oi_1 _10731_ (.A1(_05761_),
    .A2(_05762_),
    .B1(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__a31o_1 _10732_ (.A1(_05761_),
    .A2(_05762_),
    .A3(_05781_),
    .B1(_04956_),
    .X(_05783_));
 sky130_fd_sc_hd__or2_1 _10733_ (.A(_05782_),
    .B(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__o31ai_4 _10734_ (.A1(_05485_),
    .A2(_05759_),
    .A3(_05760_),
    .B1(_05784_),
    .Y(net159));
 sky130_fd_sc_hd__nand2_1 _10735_ (.A(net125),
    .B(_05760_),
    .Y(_05785_));
 sky130_fd_sc_hd__or2_1 _10736_ (.A(net125),
    .B(_05760_),
    .X(_05786_));
 sky130_fd_sc_hd__inv_2 _10737_ (.A(_05761_),
    .Y(_05787_));
 sky130_fd_sc_hd__o21ai_1 _10738_ (.A1(_05752_),
    .A2(_05787_),
    .B1(_05780_),
    .Y(_05788_));
 sky130_fd_sc_hd__o21ai_1 _10739_ (.A1(_05752_),
    .A2(_05780_),
    .B1(_05756_),
    .Y(_05789_));
 sky130_fd_sc_hd__or2_1 _10740_ (.A(net53),
    .B(net21),
    .X(_05790_));
 sky130_fd_sc_hd__nand2_1 _10741_ (.A(net53),
    .B(net21),
    .Y(_05791_));
 sky130_fd_sc_hd__nand2_1 _10742_ (.A(_05790_),
    .B(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__xor2_1 _10743_ (.A(net80),
    .B(net77),
    .X(_05793_));
 sky130_fd_sc_hd__nor2_1 _10744_ (.A(_04773_),
    .B(_05793_),
    .Y(_05794_));
 sky130_fd_sc_hd__o21a_1 _10745_ (.A1(_04759_),
    .A2(_04773_),
    .B1(_05793_),
    .X(_05795_));
 sky130_fd_sc_hd__a21oi_1 _10746_ (.A1(net79),
    .A2(_05794_),
    .B1(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hd__and3b_1 _10747_ (.A_N(_05796_),
    .B(net78),
    .C(_05768_),
    .X(_05797_));
 sky130_fd_sc_hd__a21boi_1 _10748_ (.A1(net78),
    .A2(_05768_),
    .B1_N(_05796_),
    .Y(_05798_));
 sky130_fd_sc_hd__or2_1 _10749_ (.A(_05797_),
    .B(_05798_),
    .X(_05799_));
 sky130_fd_sc_hd__a21oi_1 _10750_ (.A1(_05770_),
    .A2(_05773_),
    .B1(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hd__and3_1 _10751_ (.A(_05770_),
    .B(_05773_),
    .C(_05799_),
    .X(_05801_));
 sky130_fd_sc_hd__nor2_1 _10752_ (.A(_05800_),
    .B(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__xor2_1 _10753_ (.A(_05792_),
    .B(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__a21boi_1 _10754_ (.A1(_05763_),
    .A2(_05775_),
    .B1_N(_05764_),
    .Y(_05804_));
 sky130_fd_sc_hd__nor2_1 _10755_ (.A(_05803_),
    .B(_05804_),
    .Y(_05805_));
 sky130_fd_sc_hd__nand2_1 _10756_ (.A(_05803_),
    .B(_05804_),
    .Y(_05806_));
 sky130_fd_sc_hd__and2b_1 _10757_ (.A_N(_05805_),
    .B(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__xnor2_1 _10758_ (.A(_05778_),
    .B(_05807_),
    .Y(_05808_));
 sky130_fd_sc_hd__a21o_1 _10759_ (.A1(_05788_),
    .A2(_05789_),
    .B1(_05808_),
    .X(_05809_));
 sky130_fd_sc_hd__a31oi_1 _10760_ (.A1(_05808_),
    .A2(_05788_),
    .A3(_05789_),
    .B1(_04956_),
    .Y(_05810_));
 sky130_fd_sc_hd__a32o_1 _10761_ (.A1(_04464_),
    .A2(_05785_),
    .A3(_05786_),
    .B1(_05809_),
    .B2(_05810_),
    .X(net160));
 sky130_fd_sc_hd__nand2_1 _10762_ (.A(_05778_),
    .B(_05807_),
    .Y(_05811_));
 sky130_fd_sc_hd__and2_1 _10763_ (.A(net81),
    .B(_05738_),
    .X(_05812_));
 sky130_fd_sc_hd__nor2_1 _10764_ (.A(net81),
    .B(_05738_),
    .Y(_05813_));
 sky130_fd_sc_hd__or2_1 _10765_ (.A(_05812_),
    .B(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__nor2_1 _10766_ (.A(net77),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__inv_2 _10767_ (.A(net80),
    .Y(_05816_));
 sky130_fd_sc_hd__o21a_1 _10768_ (.A1(_05816_),
    .A2(net77),
    .B1(_05814_),
    .X(_05817_));
 sky130_fd_sc_hd__a21oi_1 _10769_ (.A1(net80),
    .A2(_05815_),
    .B1(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__or3_1 _10770_ (.A(_04759_),
    .B(_05794_),
    .C(_05818_),
    .X(_05819_));
 sky130_fd_sc_hd__o21ai_1 _10771_ (.A1(_04759_),
    .A2(_05794_),
    .B1(_05818_),
    .Y(_05820_));
 sky130_fd_sc_hd__nand2_1 _10772_ (.A(_05819_),
    .B(_05820_),
    .Y(_05821_));
 sky130_fd_sc_hd__o21bai_1 _10773_ (.A1(_05797_),
    .A2(_05800_),
    .B1_N(_05821_),
    .Y(_05822_));
 sky130_fd_sc_hd__or3b_1 _10774_ (.A(_05797_),
    .B(_05800_),
    .C_N(_05821_),
    .X(_05823_));
 sky130_fd_sc_hd__and2_1 _10775_ (.A(_05822_),
    .B(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__nor2_1 _10776_ (.A(net54),
    .B(net22),
    .Y(_05825_));
 sky130_fd_sc_hd__and2_1 _10777_ (.A(net54),
    .B(net22),
    .X(_05826_));
 sky130_fd_sc_hd__nor2_1 _10778_ (.A(_05825_),
    .B(_05826_),
    .Y(_05827_));
 sky130_fd_sc_hd__xnor2_1 _10779_ (.A(_05824_),
    .B(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__a21bo_1 _10780_ (.A1(_05790_),
    .A2(_05802_),
    .B1_N(_05791_),
    .X(_05829_));
 sky130_fd_sc_hd__xnor2_1 _10781_ (.A(_05828_),
    .B(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__nand2_1 _10782_ (.A(_05805_),
    .B(_05830_),
    .Y(_05831_));
 sky130_fd_sc_hd__or2_1 _10783_ (.A(_05805_),
    .B(_05830_),
    .X(_05832_));
 sky130_fd_sc_hd__nand2_1 _10784_ (.A(_05831_),
    .B(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__nand3_1 _10785_ (.A(_05811_),
    .B(_05809_),
    .C(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__a21o_1 _10786_ (.A1(_05811_),
    .A2(_05809_),
    .B1(_05833_),
    .X(_05835_));
 sky130_fd_sc_hd__inv_2 _10787_ (.A(net126),
    .Y(_05836_));
 sky130_fd_sc_hd__a31o_1 _10788_ (.A1(net125),
    .A2(net126),
    .A3(_05760_),
    .B1(_04687_),
    .X(_05837_));
 sky130_fd_sc_hd__a21oi_1 _10789_ (.A1(_05836_),
    .A2(_05785_),
    .B1(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__a31o_4 _10790_ (.A1(_04444_),
    .A2(_05834_),
    .A3(_05835_),
    .B1(_05838_),
    .X(net161));
 sky130_fd_sc_hd__and2b_1 _10791_ (.A_N(_05828_),
    .B(_05829_),
    .X(_05839_));
 sky130_fd_sc_hd__nand2_1 _10792_ (.A(net56),
    .B(net24),
    .Y(_05840_));
 sky130_fd_sc_hd__or2_1 _10793_ (.A(net56),
    .B(net24),
    .X(_05841_));
 sky130_fd_sc_hd__nand2_1 _10794_ (.A(_05840_),
    .B(_05841_),
    .Y(_05842_));
 sky130_fd_sc_hd__or2_1 _10795_ (.A(_05816_),
    .B(_05815_),
    .X(_05843_));
 sky130_fd_sc_hd__and2_1 _10796_ (.A(net82),
    .B(_04759_),
    .X(_05844_));
 sky130_fd_sc_hd__nor2_1 _10797_ (.A(net82),
    .B(_04759_),
    .Y(_05845_));
 sky130_fd_sc_hd__nor2_1 _10798_ (.A(_05844_),
    .B(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__and2_1 _10799_ (.A(_05738_),
    .B(_05846_),
    .X(_05847_));
 sky130_fd_sc_hd__o2bb2a_1 _10800_ (.A1_N(net81),
    .A2_N(_05847_),
    .B1(_05846_),
    .B2(_05812_),
    .X(_05848_));
 sky130_fd_sc_hd__xnor2_1 _10801_ (.A(_05843_),
    .B(_05848_),
    .Y(_05849_));
 sky130_fd_sc_hd__and3_1 _10802_ (.A(_05819_),
    .B(_05822_),
    .C(_05849_),
    .X(_05850_));
 sky130_fd_sc_hd__a21o_1 _10803_ (.A1(_05819_),
    .A2(_05822_),
    .B1(_05849_),
    .X(_05851_));
 sky130_fd_sc_hd__and2b_1 _10804_ (.A_N(_05850_),
    .B(_05851_),
    .X(_05852_));
 sky130_fd_sc_hd__xor2_1 _10805_ (.A(_05842_),
    .B(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__a21oi_1 _10806_ (.A1(_05824_),
    .A2(_05827_),
    .B1(_05826_),
    .Y(_05854_));
 sky130_fd_sc_hd__xor2_1 _10807_ (.A(_05853_),
    .B(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__and2_1 _10808_ (.A(_05839_),
    .B(_05855_),
    .X(_05856_));
 sky130_fd_sc_hd__nor2_1 _10809_ (.A(_05839_),
    .B(_05855_),
    .Y(_05857_));
 sky130_fd_sc_hd__or2_1 _10810_ (.A(_05856_),
    .B(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__a21oi_2 _10811_ (.A1(_05831_),
    .A2(_05835_),
    .B1(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__a31o_1 _10812_ (.A1(_05831_),
    .A2(_05835_),
    .A3(_05858_),
    .B1(_04956_),
    .X(_05860_));
 sky130_fd_sc_hd__and4_1 _10813_ (.A(net125),
    .B(net126),
    .C(net128),
    .D(_05760_),
    .X(_05861_));
 sky130_fd_sc_hd__a31o_1 _10814_ (.A1(net125),
    .A2(net126),
    .A3(_05760_),
    .B1(net128),
    .X(_05862_));
 sky130_fd_sc_hd__or3b_2 _10815_ (.A(_04688_),
    .B(_05861_),
    .C_N(_05862_),
    .X(_05863_));
 sky130_fd_sc_hd__o21ai_4 _10816_ (.A1(_05859_),
    .A2(_05860_),
    .B1(_05863_),
    .Y(net163));
 sky130_fd_sc_hd__a21bo_1 _10817_ (.A1(_05841_),
    .A2(_05852_),
    .B1_N(_05840_),
    .X(_05864_));
 sky130_fd_sc_hd__o21a_1 _10818_ (.A1(_05843_),
    .A2(_05848_),
    .B1(_05851_),
    .X(_05865_));
 sky130_fd_sc_hd__xor2_1 _10819_ (.A(_05864_),
    .B(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__xor2_2 _10820_ (.A(net83),
    .B(net80),
    .X(_05867_));
 sky130_fd_sc_hd__xnor2_1 _10821_ (.A(_05866_),
    .B(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__nor2_1 _10822_ (.A(_05844_),
    .B(_05847_),
    .Y(_05869_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(_05844_),
    .A1(_05869_),
    .S(net81),
    .X(_05870_));
 sky130_fd_sc_hd__xnor2_1 _10824_ (.A(_05868_),
    .B(_05870_),
    .Y(_05871_));
 sky130_fd_sc_hd__nor2_1 _10825_ (.A(_05853_),
    .B(_05854_),
    .Y(_05872_));
 sky130_fd_sc_hd__xnor2_4 _10826_ (.A(net57),
    .B(net25),
    .Y(_05873_));
 sky130_fd_sc_hd__xnor2_1 _10827_ (.A(_05872_),
    .B(_05873_),
    .Y(_05874_));
 sky130_fd_sc_hd__xnor2_1 _10828_ (.A(_05871_),
    .B(_05874_),
    .Y(_05875_));
 sky130_fd_sc_hd__o21ai_1 _10829_ (.A1(_05856_),
    .A2(_05859_),
    .B1(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__o31a_1 _10830_ (.A1(_05856_),
    .A2(_05859_),
    .A3(_05875_),
    .B1(_04443_),
    .X(_05877_));
 sky130_fd_sc_hd__xor2_1 _10831_ (.A(net129),
    .B(_05861_),
    .X(_05878_));
 sky130_fd_sc_hd__a22o_4 _10832_ (.A1(_05876_),
    .A2(_05877_),
    .B1(_05878_),
    .B2(_04464_),
    .X(net164));
 sky130_fd_sc_hd__o21ba_1 _10833_ (.A1(_04449_),
    .A2(net1786),
    .B1_N(net138),
    .X(_00000_));
 sky130_fd_sc_hd__or3_1 _10834_ (.A(\cand_x[2] ),
    .B(\cand_x[1] ),
    .C(\cand_x[0] ),
    .X(_05879_));
 sky130_fd_sc_hd__inv_2 _10835_ (.A(_04475_),
    .Y(_05880_));
 sky130_fd_sc_hd__o31a_1 _10836_ (.A1(\cand_x[4] ),
    .A2(\cand_x[3] ),
    .A3(_05879_),
    .B1(_05880_),
    .X(_05881_));
 sky130_fd_sc_hd__or4_1 _10837_ (.A(\cand_y[3] ),
    .B(\cand_y[2] ),
    .C(\cand_y[1] ),
    .D(\cand_y[0] ),
    .X(_05882_));
 sky130_fd_sc_hd__o211ai_1 _10838_ (.A1(\cand_y[4] ),
    .A2(_05882_),
    .B1(_04752_),
    .C1(\cand_y[5] ),
    .Y(_05883_));
 sky130_fd_sc_hd__o221a_1 _10839_ (.A1(\cand_x[5] ),
    .A2(_05880_),
    .B1(\cand_y[5] ),
    .B2(_04752_),
    .C1(_05883_),
    .X(_05884_));
 sky130_fd_sc_hd__a21boi_1 _10840_ (.A1(\cand_x[5] ),
    .A2(_05881_),
    .B1_N(_05884_),
    .Y(_05885_));
 sky130_fd_sc_hd__clkbuf_4 _10841_ (.A(net217),
    .X(_05886_));
 sky130_fd_sc_hd__or2_1 _10842_ (.A(_04654_),
    .B(_04459_),
    .X(_05887_));
 sky130_fd_sc_hd__or2b_1 _10843_ (.A(_04670_),
    .B_N(_04692_),
    .X(_05888_));
 sky130_fd_sc_hd__nor4b_1 _10844_ (.A(_04653_),
    .B(_04458_),
    .C(_04691_),
    .D_N(_04669_),
    .Y(_05889_));
 sky130_fd_sc_hd__buf_12 _10845_ (.A(net260),
    .X(_05890_));
 sky130_fd_sc_hd__and4bb_2 _10846_ (.A_N(_04420_),
    .B_N(\pixel_cnt[2] ),
    .C(\pixel_cnt[3] ),
    .D(_04421_),
    .X(_05891_));
 sky130_fd_sc_hd__clkbuf_16 _10847_ (.A(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__clkbuf_16 _10848_ (.A(_05892_),
    .X(_05893_));
 sky130_fd_sc_hd__nor4b_1 _10849_ (.A(_04653_),
    .B(_04458_),
    .C(_04669_),
    .D_N(_04691_),
    .Y(_05894_));
 sky130_fd_sc_hd__buf_12 _10850_ (.A(net258),
    .X(_05895_));
 sky130_fd_sc_hd__buf_8 _10851_ (.A(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__a2111o_2 _10852_ (.A1(_05887_),
    .A2(_05888_),
    .B1(_05890_),
    .C1(_05893_),
    .D1(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__and2_1 _10853_ (.A(_04654_),
    .B(_04459_),
    .X(_05898_));
 sky130_fd_sc_hd__or4_4 _10854_ (.A(_04425_),
    .B(_04426_),
    .C(_04427_),
    .D(_04428_),
    .X(_05899_));
 sky130_fd_sc_hd__and4bb_4 _10855_ (.A_N(_04420_),
    .B_N(_04421_),
    .C(\pixel_cnt[2] ),
    .D(\pixel_cnt[3] ),
    .X(_05900_));
 sky130_fd_sc_hd__buf_12 _10856_ (.A(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__buf_12 _10857_ (.A(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__and4bb_2 _10858_ (.A_N(_04421_),
    .B_N(\pixel_cnt[2] ),
    .C(\pixel_cnt[3] ),
    .D(_04420_),
    .X(_05903_));
 sky130_fd_sc_hd__buf_8 _10859_ (.A(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__buf_12 _10860_ (.A(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__or4_4 _10861_ (.A(_05898_),
    .B(_05899_),
    .C(_05902_),
    .D(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__or2_2 _10862_ (.A(_05897_),
    .B(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__clkbuf_8 _10863_ (.A(_05907_),
    .X(_05908_));
 sky130_fd_sc_hd__buf_12 _10864_ (.A(_05891_),
    .X(_05909_));
 sky130_fd_sc_hd__buf_12 _10865_ (.A(_05909_),
    .X(_05910_));
 sky130_fd_sc_hd__clkbuf_16 _10866_ (.A(_05910_),
    .X(_05911_));
 sky130_fd_sc_hd__buf_6 _10867_ (.A(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__and4bb_4 _10868_ (.A_N(_04426_),
    .B_N(_04427_),
    .C(_04428_),
    .D(_04425_),
    .X(_05913_));
 sky130_fd_sc_hd__buf_4 _10869_ (.A(net253),
    .X(_05914_));
 sky130_fd_sc_hd__clkbuf_8 _10870_ (.A(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__buf_6 _10871_ (.A(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__and4b_4 _10872_ (.A_N(_04669_),
    .B(_04691_),
    .C(_04653_),
    .D(_04458_),
    .X(_05917_));
 sky130_fd_sc_hd__clkbuf_8 _10873_ (.A(_05917_),
    .X(_05918_));
 sky130_fd_sc_hd__clkbuf_16 _10874_ (.A(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__and4bb_4 _10875_ (.A_N(_05053_),
    .B_N(_05052_),
    .C(_05051_),
    .D(_05054_),
    .X(_05920_));
 sky130_fd_sc_hd__buf_6 _10876_ (.A(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__buf_12 _10877_ (.A(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__buf_8 _10878_ (.A(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__and3_1 _10879_ (.A(\cur_mb_mem[171][7] ),
    .B(_05919_),
    .C(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__buf_4 _10880_ (.A(_05915_),
    .X(_05925_));
 sky130_fd_sc_hd__nor4_4 _10881_ (.A(_04425_),
    .B(_04426_),
    .C(_04427_),
    .D(_04428_),
    .Y(_05926_));
 sky130_fd_sc_hd__and2_1 _10882_ (.A(net250),
    .B(_05900_),
    .X(_05927_));
 sky130_fd_sc_hd__buf_6 _10883_ (.A(_05927_),
    .X(_05928_));
 sky130_fd_sc_hd__a32o_1 _10884_ (.A1(\cur_mb_mem[88][7] ),
    .A2(_05896_),
    .A3(_05925_),
    .B1(_05928_),
    .B2(\cur_mb_mem[12][7] ),
    .X(_05929_));
 sky130_fd_sc_hd__a311o_1 _10885_ (.A1(\cur_mb_mem[89][7] ),
    .A2(_05912_),
    .A3(_05916_),
    .B1(_05924_),
    .C1(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__clkbuf_16 _10886_ (.A(_05904_),
    .X(_05931_));
 sky130_fd_sc_hd__nor4b_1 _10887_ (.A(_05053_),
    .B(_05054_),
    .C(_05052_),
    .D_N(_05051_),
    .Y(_05932_));
 sky130_fd_sc_hd__clkbuf_16 _10888_ (.A(net245),
    .X(_05933_));
 sky130_fd_sc_hd__and2_4 _10889_ (.A(_05931_),
    .B(_05933_),
    .X(_05934_));
 sky130_fd_sc_hd__clkbuf_16 _10890_ (.A(net247),
    .X(_05935_));
 sky130_fd_sc_hd__and2_2 _10891_ (.A(_05910_),
    .B(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__buf_12 _10892_ (.A(_05901_),
    .X(_05937_));
 sky130_fd_sc_hd__buf_8 _10893_ (.A(_05937_),
    .X(_05938_));
 sky130_fd_sc_hd__and4b_4 _10894_ (.A_N(_05054_),
    .B(\pixel_cnt[7] ),
    .C(\pixel_cnt[6] ),
    .D(\pixel_cnt[4] ),
    .X(_05939_));
 sky130_fd_sc_hd__clkbuf_4 _10895_ (.A(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__buf_8 _10896_ (.A(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__clkbuf_8 _10897_ (.A(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__and4b_4 _10898_ (.A_N(_04420_),
    .B(_04421_),
    .C(\pixel_cnt[2] ),
    .D(\pixel_cnt[3] ),
    .X(_05943_));
 sky130_fd_sc_hd__buf_6 _10899_ (.A(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__buf_8 _10900_ (.A(_05944_),
    .X(_05945_));
 sky130_fd_sc_hd__buf_8 _10901_ (.A(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__clkbuf_8 _10902_ (.A(_05940_),
    .X(_05947_));
 sky130_fd_sc_hd__buf_6 _10903_ (.A(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__and3_1 _10904_ (.A(\cur_mb_mem[221][7] ),
    .B(_05946_),
    .C(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__a31o_2 _10905_ (.A1(\cur_mb_mem[220][7] ),
    .A2(_05938_),
    .A3(_05942_),
    .B1(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__a221o_1 _10906_ (.A1(\cur_mb_mem[138][7] ),
    .A2(_05934_),
    .B1(_05936_),
    .B2(\cur_mb_mem[137][7] ),
    .C1(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__and4b_4 _10907_ (.A_N(_04421_),
    .B(\pixel_cnt[2] ),
    .C(\pixel_cnt[3] ),
    .D(_04420_),
    .X(_05952_));
 sky130_fd_sc_hd__buf_4 _10908_ (.A(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__buf_8 _10909_ (.A(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__buf_4 _10910_ (.A(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__clkbuf_8 _10911_ (.A(_05923_),
    .X(_05956_));
 sky130_fd_sc_hd__buf_12 _10912_ (.A(_05904_),
    .X(_05957_));
 sky130_fd_sc_hd__buf_8 _10913_ (.A(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__buf_6 _10914_ (.A(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__and3_1 _10915_ (.A(\cur_mb_mem[90][7] ),
    .B(_05959_),
    .C(_05925_),
    .X(_05960_));
 sky130_fd_sc_hd__buf_8 _10916_ (.A(_05946_),
    .X(_05961_));
 sky130_fd_sc_hd__or4b_1 _10917_ (.A(_04653_),
    .B(_04669_),
    .C(_04691_),
    .D_N(_04458_),
    .X(_05962_));
 sky130_fd_sc_hd__buf_8 _10918_ (.A(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__or4b_1 _10919_ (.A(_04425_),
    .B(_04426_),
    .C(_04428_),
    .D_N(_04427_),
    .X(_05964_));
 sky130_fd_sc_hd__buf_8 _10920_ (.A(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__nor2_8 _10921_ (.A(_05963_),
    .B(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__a32o_1 _10922_ (.A1(\cur_mb_mem[93][7] ),
    .A2(_05925_),
    .A3(_05961_),
    .B1(_05966_),
    .B2(\cur_mb_mem[129][7] ),
    .X(_05967_));
 sky130_fd_sc_hd__a311o_1 _10923_ (.A1(\cur_mb_mem[174][7] ),
    .A2(_05955_),
    .A3(_05956_),
    .B1(_05960_),
    .C1(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__nor4_1 _10924_ (.A(_04653_),
    .B(_04458_),
    .C(_04669_),
    .D(_04691_),
    .Y(_05969_));
 sky130_fd_sc_hd__buf_12 _10925_ (.A(net241),
    .X(_05970_));
 sky130_fd_sc_hd__buf_6 _10926_ (.A(_05970_),
    .X(_05971_));
 sky130_fd_sc_hd__buf_6 _10927_ (.A(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__buf_8 _10928_ (.A(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__nor4b_1 _10929_ (.A(_04426_),
    .B(_04427_),
    .C(_04428_),
    .D_N(_04425_),
    .Y(_05974_));
 sky130_fd_sc_hd__buf_8 _10930_ (.A(net234),
    .X(_05975_));
 sky130_fd_sc_hd__buf_12 _10931_ (.A(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__and4bb_4 _10932_ (.A_N(_04426_),
    .B_N(_04428_),
    .C(_05051_),
    .D(_04425_),
    .X(_05977_));
 sky130_fd_sc_hd__buf_8 _10933_ (.A(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__buf_8 _10934_ (.A(_05978_),
    .X(_05979_));
 sky130_fd_sc_hd__clkbuf_8 _10935_ (.A(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__and3_1 _10936_ (.A(\cur_mb_mem[156][7] ),
    .B(_05938_),
    .C(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__buf_12 _10937_ (.A(net257),
    .X(_05982_));
 sky130_fd_sc_hd__and4bb_4 _10938_ (.A_N(_05053_),
    .B_N(_05051_),
    .C(_05052_),
    .D(_05054_),
    .X(_05983_));
 sky130_fd_sc_hd__buf_4 _10939_ (.A(_05983_),
    .X(_05984_));
 sky130_fd_sc_hd__and2_4 _10940_ (.A(_05982_),
    .B(_05984_),
    .X(_05985_));
 sky130_fd_sc_hd__a32o_2 _10941_ (.A1(\cur_mb_mem[154][7] ),
    .A2(_05959_),
    .A3(_05980_),
    .B1(_05985_),
    .B2(\cur_mb_mem[104][7] ),
    .X(_05986_));
 sky130_fd_sc_hd__a311o_1 _10942_ (.A1(\cur_mb_mem[16][7] ),
    .A2(_05973_),
    .A3(_05976_),
    .B1(_05981_),
    .C1(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__or4_1 _10943_ (.A(_05930_),
    .B(_05951_),
    .C(_05968_),
    .D(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__clkbuf_8 _10944_ (.A(_05938_),
    .X(_05989_));
 sky130_fd_sc_hd__nor2_8 _10945_ (.A(_05899_),
    .B(_05963_),
    .Y(_05990_));
 sky130_fd_sc_hd__a32o_1 _10946_ (.A1(\cur_mb_mem[172][7] ),
    .A2(_05989_),
    .A3(_05956_),
    .B1(_05990_),
    .B2(\cur_mb_mem[1][7] ),
    .X(_05991_));
 sky130_fd_sc_hd__nor4b_1 _10947_ (.A(_04653_),
    .B(_04669_),
    .C(_04691_),
    .D_N(_04458_),
    .Y(_05992_));
 sky130_fd_sc_hd__clkbuf_16 _10948_ (.A(net229),
    .X(_05993_));
 sky130_fd_sc_hd__clkbuf_16 _10949_ (.A(_05993_),
    .X(_05994_));
 sky130_fd_sc_hd__buf_12 _10950_ (.A(net229),
    .X(_05995_));
 sky130_fd_sc_hd__and4b_2 _10951_ (.A_N(_05053_),
    .B(\pixel_cnt[5] ),
    .C(_05051_),
    .D(_05052_),
    .X(_05996_));
 sky130_fd_sc_hd__buf_4 _10952_ (.A(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__and2_4 _10953_ (.A(_05995_),
    .B(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__a32o_1 _10954_ (.A1(\cur_mb_mem[49][7] ),
    .A2(_05058_),
    .A3(_05994_),
    .B1(_05998_),
    .B2(\cur_mb_mem[225][7] ),
    .X(_05999_));
 sky130_fd_sc_hd__buf_12 _10955_ (.A(_05953_),
    .X(_06000_));
 sky130_fd_sc_hd__buf_12 _10956_ (.A(net235),
    .X(_06001_));
 sky130_fd_sc_hd__and2_4 _10957_ (.A(_06000_),
    .B(_06001_),
    .X(_06002_));
 sky130_fd_sc_hd__buf_6 _10958_ (.A(_05917_),
    .X(_06003_));
 sky130_fd_sc_hd__nor4b_1 _10959_ (.A(_05053_),
    .B(_04427_),
    .C(_05052_),
    .D_N(_05054_),
    .Y(_06004_));
 sky130_fd_sc_hd__clkbuf_8 _10960_ (.A(net225),
    .X(_06005_));
 sky130_fd_sc_hd__and2_4 _10961_ (.A(_06003_),
    .B(_06005_),
    .X(_06006_));
 sky130_fd_sc_hd__a22o_2 _10962_ (.A1(\cur_mb_mem[30][7] ),
    .A2(_06002_),
    .B1(_06006_),
    .B2(\cur_mb_mem[43][7] ),
    .X(_06007_));
 sky130_fd_sc_hd__clkbuf_8 _10963_ (.A(net253),
    .X(_06008_));
 sky130_fd_sc_hd__buf_12 _10964_ (.A(net240),
    .X(_06009_));
 sky130_fd_sc_hd__and2_4 _10965_ (.A(_06008_),
    .B(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__clkbuf_16 _10966_ (.A(_05944_),
    .X(_06011_));
 sky130_fd_sc_hd__and4b_1 _10967_ (.A_N(_05052_),
    .B(_05051_),
    .C(_05054_),
    .D(_05053_),
    .X(_06012_));
 sky130_fd_sc_hd__buf_6 _10968_ (.A(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__and2_2 _10969_ (.A(_06011_),
    .B(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__a22o_1 _10970_ (.A1(\cur_mb_mem[80][7] ),
    .A2(_06010_),
    .B1(_06014_),
    .B2(\cur_mb_mem[189][7] ),
    .X(_06015_));
 sky130_fd_sc_hd__or4_1 _10971_ (.A(_05991_),
    .B(_05999_),
    .C(_06007_),
    .D(_06015_),
    .X(_06016_));
 sky130_fd_sc_hd__and2_4 _10972_ (.A(_05937_),
    .B(_05975_),
    .X(_06017_));
 sky130_fd_sc_hd__buf_6 _10973_ (.A(_06012_),
    .X(_06018_));
 sky130_fd_sc_hd__buf_6 _10974_ (.A(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__and2_4 _10975_ (.A(_06019_),
    .B(_05995_),
    .X(_06020_));
 sky130_fd_sc_hd__nor4b_1 _10976_ (.A(_05053_),
    .B(_05054_),
    .C(_05051_),
    .D_N(_05052_),
    .Y(_06021_));
 sky130_fd_sc_hd__buf_4 _10977_ (.A(net224),
    .X(_06022_));
 sky130_fd_sc_hd__clkbuf_8 _10978_ (.A(_06022_),
    .X(_06023_));
 sky130_fd_sc_hd__buf_8 _10979_ (.A(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__buf_8 _10980_ (.A(_05955_),
    .X(_06025_));
 sky130_fd_sc_hd__buf_12 _10981_ (.A(net262),
    .X(_06026_));
 sky130_fd_sc_hd__buf_4 _10982_ (.A(_05983_),
    .X(_06027_));
 sky130_fd_sc_hd__and2_4 _10983_ (.A(_06026_),
    .B(_06027_),
    .X(_06028_));
 sky130_fd_sc_hd__a32o_1 _10984_ (.A1(\cur_mb_mem[78][7] ),
    .A2(_06024_),
    .A3(_06025_),
    .B1(_06028_),
    .B2(\cur_mb_mem[100][7] ),
    .X(_06029_));
 sky130_fd_sc_hd__a221o_1 _10985_ (.A1(\cur_mb_mem[28][7] ),
    .A2(_06017_),
    .B1(_06020_),
    .B2(\cur_mb_mem[177][7] ),
    .C1(_06029_),
    .X(_06030_));
 sky130_fd_sc_hd__and2_4 _10986_ (.A(_05909_),
    .B(_06005_),
    .X(_06031_));
 sky130_fd_sc_hd__buf_8 _10987_ (.A(_04429_),
    .X(_06032_));
 sky130_fd_sc_hd__buf_6 _10988_ (.A(_05943_),
    .X(_06033_));
 sky130_fd_sc_hd__and2_4 _10989_ (.A(_06032_),
    .B(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__clkbuf_8 _10990_ (.A(_05959_),
    .X(_06035_));
 sky130_fd_sc_hd__buf_8 _10991_ (.A(_06018_),
    .X(_06036_));
 sky130_fd_sc_hd__buf_4 _10992_ (.A(_06036_),
    .X(_06037_));
 sky130_fd_sc_hd__buf_12 _10993_ (.A(_05892_),
    .X(_06038_));
 sky130_fd_sc_hd__buf_8 _10994_ (.A(_06018_),
    .X(_06039_));
 sky130_fd_sc_hd__and2_4 _10995_ (.A(_06038_),
    .B(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__a32o_1 _10996_ (.A1(\cur_mb_mem[186][7] ),
    .A2(_06035_),
    .A3(_06037_),
    .B1(_06040_),
    .B2(\cur_mb_mem[185][7] ),
    .X(_06041_));
 sky130_fd_sc_hd__a221o_2 _10997_ (.A1(\cur_mb_mem[41][7] ),
    .A2(_06031_),
    .B1(_06034_),
    .B2(\cur_mb_mem[253][7] ),
    .C1(_06041_),
    .X(_06042_));
 sky130_fd_sc_hd__or4_1 _10998_ (.A(_05988_),
    .B(_06016_),
    .C(_06030_),
    .D(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__buf_8 _10999_ (.A(net226),
    .X(_06044_));
 sky130_fd_sc_hd__buf_4 _11000_ (.A(_05983_),
    .X(_06045_));
 sky130_fd_sc_hd__clkbuf_16 _11001_ (.A(_05952_),
    .X(_06046_));
 sky130_fd_sc_hd__and2_4 _11002_ (.A(_06045_),
    .B(_06046_),
    .X(_06047_));
 sky130_fd_sc_hd__a32o_1 _11003_ (.A1(\cur_mb_mem[32][7] ),
    .A2(_06044_),
    .A3(_05973_),
    .B1(_06047_),
    .B2(\cur_mb_mem[110][7] ),
    .X(_06048_));
 sky130_fd_sc_hd__buf_8 _11004_ (.A(_05919_),
    .X(_06049_));
 sky130_fd_sc_hd__and4b_4 _11005_ (.A_N(_05051_),
    .B(_05052_),
    .C(_05053_),
    .D(_05054_),
    .X(_06050_));
 sky130_fd_sc_hd__buf_4 _11006_ (.A(_06050_),
    .X(_06051_));
 sky130_fd_sc_hd__clkbuf_8 _11007_ (.A(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__clkbuf_8 _11008_ (.A(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__and3_2 _11009_ (.A(\cur_mb_mem[122][7] ),
    .B(_05959_),
    .C(_06053_),
    .X(_06054_));
 sky130_fd_sc_hd__a31o_2 _11010_ (.A1(\cur_mb_mem[251][7] ),
    .A2(_04432_),
    .A3(_06049_),
    .B1(_06054_),
    .X(_06055_));
 sky130_fd_sc_hd__buf_8 _11011_ (.A(_05944_),
    .X(_06056_));
 sky130_fd_sc_hd__buf_6 _11012_ (.A(_06022_),
    .X(_06057_));
 sky130_fd_sc_hd__and2_4 _11013_ (.A(_06056_),
    .B(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__a32o_1 _11014_ (.A1(\cur_mb_mem[48][7] ),
    .A2(_05058_),
    .A3(_05973_),
    .B1(_06058_),
    .B2(\cur_mb_mem[77][7] ),
    .X(_06059_));
 sky130_fd_sc_hd__and4bb_4 _11015_ (.A_N(\pixel_cnt[2] ),
    .B_N(\pixel_cnt[3] ),
    .C(_04420_),
    .D(_04421_),
    .X(_06060_));
 sky130_fd_sc_hd__buf_12 _11016_ (.A(_06060_),
    .X(_06061_));
 sky130_fd_sc_hd__buf_8 _11017_ (.A(_06061_),
    .X(_06062_));
 sky130_fd_sc_hd__buf_12 _11018_ (.A(_06062_),
    .X(_06063_));
 sky130_fd_sc_hd__buf_8 _11019_ (.A(_06063_),
    .X(_06064_));
 sky130_fd_sc_hd__buf_4 _11020_ (.A(_05997_),
    .X(_06065_));
 sky130_fd_sc_hd__buf_4 _11021_ (.A(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__buf_4 _11022_ (.A(_06066_),
    .X(_06067_));
 sky130_fd_sc_hd__clkbuf_16 _11023_ (.A(_04422_),
    .X(_06068_));
 sky130_fd_sc_hd__and2_4 _11024_ (.A(_06068_),
    .B(_06027_),
    .X(_06069_));
 sky130_fd_sc_hd__a32o_2 _11025_ (.A1(\cur_mb_mem[227][7] ),
    .A2(_06064_),
    .A3(_06067_),
    .B1(_06069_),
    .B2(\cur_mb_mem[111][7] ),
    .X(_06070_));
 sky130_fd_sc_hd__and3_1 _11026_ (.A(\cur_mb_mem[92][7] ),
    .B(_05989_),
    .C(_05925_),
    .X(_06071_));
 sky130_fd_sc_hd__a31o_1 _11027_ (.A1(\cur_mb_mem[57][7] ),
    .A2(_05058_),
    .A3(_05912_),
    .B1(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__or4_1 _11028_ (.A(_06055_),
    .B(_06059_),
    .C(_06070_),
    .D(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__buf_12 _11029_ (.A(net243),
    .X(_06074_));
 sky130_fd_sc_hd__and2_2 _11030_ (.A(_06074_),
    .B(_05933_),
    .X(_06075_));
 sky130_fd_sc_hd__clkbuf_16 _11031_ (.A(net228),
    .X(_06076_));
 sky130_fd_sc_hd__and2_4 _11032_ (.A(_06027_),
    .B(_06076_),
    .X(_06077_));
 sky130_fd_sc_hd__nor4b_2 _11033_ (.A(_04458_),
    .B(_04669_),
    .C(_04691_),
    .D_N(_04420_),
    .Y(_06078_));
 sky130_fd_sc_hd__buf_12 _11034_ (.A(net223),
    .X(_06079_));
 sky130_fd_sc_hd__clkbuf_16 _11035_ (.A(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__and4bb_4 _11036_ (.A_N(_05053_),
    .B_N(_05054_),
    .C(_05051_),
    .D(_05052_),
    .X(_06081_));
 sky130_fd_sc_hd__clkbuf_16 _11037_ (.A(_06081_),
    .X(_06082_));
 sky130_fd_sc_hd__and2_4 _11038_ (.A(_06080_),
    .B(_06082_),
    .X(_06083_));
 sky130_fd_sc_hd__a32o_1 _11039_ (.A1(\cur_mb_mem[240][7] ),
    .A2(_04432_),
    .A3(_05973_),
    .B1(_06083_),
    .B2(\cur_mb_mem[194][7] ),
    .X(_06084_));
 sky130_fd_sc_hd__a221o_1 _11040_ (.A1(\cur_mb_mem[128][7] ),
    .A2(_06075_),
    .B1(_06077_),
    .B2(\cur_mb_mem[97][7] ),
    .C1(_06084_),
    .X(_06085_));
 sky130_fd_sc_hd__buf_12 _11041_ (.A(_06061_),
    .X(_06086_));
 sky130_fd_sc_hd__buf_8 _11042_ (.A(_06005_),
    .X(_06087_));
 sky130_fd_sc_hd__and2_4 _11043_ (.A(_06086_),
    .B(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__a32o_1 _11044_ (.A1(\cur_mb_mem[94][7] ),
    .A2(_05916_),
    .A3(_06025_),
    .B1(_06088_),
    .B2(\cur_mb_mem[35][7] ),
    .X(_06089_));
 sky130_fd_sc_hd__or4_1 _11045_ (.A(_06048_),
    .B(_06073_),
    .C(_06085_),
    .D(_06089_),
    .X(_06090_));
 sky130_fd_sc_hd__buf_6 _11046_ (.A(_06081_),
    .X(_06091_));
 sky130_fd_sc_hd__buf_6 _11047_ (.A(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__buf_6 _11048_ (.A(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__buf_6 _11049_ (.A(_06093_),
    .X(_06094_));
 sky130_fd_sc_hd__and4b_4 _11050_ (.A_N(_04691_),
    .B(\pixel_cnt[2] ),
    .C(_04421_),
    .D(_04420_),
    .X(_06095_));
 sky130_fd_sc_hd__buf_6 _11051_ (.A(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__buf_4 _11052_ (.A(_06096_),
    .X(_06097_));
 sky130_fd_sc_hd__buf_4 _11053_ (.A(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__buf_8 _11054_ (.A(_04422_),
    .X(_06099_));
 sky130_fd_sc_hd__and2_1 _11055_ (.A(_06099_),
    .B(_06050_),
    .X(_06100_));
 sky130_fd_sc_hd__clkbuf_8 _11056_ (.A(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__a32o_1 _11057_ (.A1(\cur_mb_mem[199][7] ),
    .A2(_06094_),
    .A3(_06098_),
    .B1(_06101_),
    .B2(\cur_mb_mem[127][7] ),
    .X(_06102_));
 sky130_fd_sc_hd__buf_4 _11058_ (.A(_06098_),
    .X(_06103_));
 sky130_fd_sc_hd__and3_1 _11059_ (.A(\cur_mb_mem[236][7] ),
    .B(_05938_),
    .C(_06066_),
    .X(_06104_));
 sky130_fd_sc_hd__a31o_1 _11060_ (.A1(\cur_mb_mem[183][7] ),
    .A2(_06037_),
    .A3(_06103_),
    .B1(_06104_),
    .X(_06105_));
 sky130_fd_sc_hd__buf_4 _11061_ (.A(_05942_),
    .X(_06106_));
 sky130_fd_sc_hd__and2_4 _11062_ (.A(_06044_),
    .B(_05954_),
    .X(_06107_));
 sky130_fd_sc_hd__a32o_1 _11063_ (.A1(\cur_mb_mem[219][7] ),
    .A2(_06049_),
    .A3(_06106_),
    .B1(_06107_),
    .B2(\cur_mb_mem[46][7] ),
    .X(_06108_));
 sky130_fd_sc_hd__and3_1 _11064_ (.A(\cur_mb_mem[238][7] ),
    .B(_05955_),
    .C(_06066_),
    .X(_06109_));
 sky130_fd_sc_hd__a31o_1 _11065_ (.A1(\cur_mb_mem[224][7] ),
    .A2(_05973_),
    .A3(_06067_),
    .B1(_06109_),
    .X(_06110_));
 sky130_fd_sc_hd__or4_1 _11066_ (.A(_06102_),
    .B(_06105_),
    .C(_06108_),
    .D(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__buf_8 _11067_ (.A(net250),
    .X(_06112_));
 sky130_fd_sc_hd__clkbuf_8 _11068_ (.A(_06112_),
    .X(_06113_));
 sky130_fd_sc_hd__and2_1 _11069_ (.A(_06113_),
    .B(_06098_),
    .X(_06114_));
 sky130_fd_sc_hd__buf_12 _11070_ (.A(_05904_),
    .X(_06115_));
 sky130_fd_sc_hd__clkbuf_4 _11071_ (.A(_05996_),
    .X(_06116_));
 sky130_fd_sc_hd__and2_4 _11072_ (.A(_06115_),
    .B(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__clkbuf_8 _11073_ (.A(_06052_),
    .X(_06118_));
 sky130_fd_sc_hd__buf_6 _11074_ (.A(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__clkbuf_16 _11075_ (.A(_06099_),
    .X(_06120_));
 sky130_fd_sc_hd__buf_6 _11076_ (.A(_06022_),
    .X(_06121_));
 sky130_fd_sc_hd__and2_4 _11077_ (.A(_06120_),
    .B(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__a32o_1 _11078_ (.A1(\cur_mb_mem[119][7] ),
    .A2(_06119_),
    .A3(_06103_),
    .B1(_06122_),
    .B2(\cur_mb_mem[79][7] ),
    .X(_06123_));
 sky130_fd_sc_hd__a221o_1 _11079_ (.A1(\cur_mb_mem[7][7] ),
    .A2(_06114_),
    .B1(_06117_),
    .B2(\cur_mb_mem[234][7] ),
    .C1(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__and2_2 _11080_ (.A(_06120_),
    .B(_05997_),
    .X(_06125_));
 sky130_fd_sc_hd__a32o_1 _11081_ (.A1(\cur_mb_mem[151][7] ),
    .A2(_05980_),
    .A3(_06103_),
    .B1(_06125_),
    .B2(\cur_mb_mem[239][7] ),
    .X(_06126_));
 sky130_fd_sc_hd__and3_1 _11082_ (.A(\cur_mb_mem[233][7] ),
    .B(_05912_),
    .C(_06067_),
    .X(_06127_));
 sky130_fd_sc_hd__a31o_1 _11083_ (.A1(\cur_mb_mem[23][7] ),
    .A2(_06103_),
    .A3(_05976_),
    .B1(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__or4_2 _11084_ (.A(_06111_),
    .B(_06124_),
    .C(_06126_),
    .D(_06128_),
    .X(_06129_));
 sky130_fd_sc_hd__and4bb_4 _11085_ (.A_N(_04653_),
    .B_N(_04691_),
    .C(_04669_),
    .D(_04421_),
    .X(_06130_));
 sky130_fd_sc_hd__buf_12 _11086_ (.A(_06130_),
    .X(_06131_));
 sky130_fd_sc_hd__buf_6 _11087_ (.A(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__clkbuf_8 _11088_ (.A(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__buf_8 _11089_ (.A(_05890_),
    .X(_06134_));
 sky130_fd_sc_hd__and2_2 _11090_ (.A(_06134_),
    .B(_05941_),
    .X(_06135_));
 sky130_fd_sc_hd__a32o_1 _11091_ (.A1(\cur_mb_mem[197][7] ),
    .A2(_06093_),
    .A3(_06133_),
    .B1(_06135_),
    .B2(\cur_mb_mem[212][7] ),
    .X(_06136_));
 sky130_fd_sc_hd__buf_8 _11092_ (.A(_05922_),
    .X(_06137_));
 sky130_fd_sc_hd__clkbuf_8 _11093_ (.A(_06050_),
    .X(_06138_));
 sky130_fd_sc_hd__and4bb_4 _11094_ (.A_N(_04421_),
    .B_N(\pixel_cnt[3] ),
    .C(\pixel_cnt[2] ),
    .D(_04420_),
    .X(_06139_));
 sky130_fd_sc_hd__buf_12 _11095_ (.A(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__and2_4 _11096_ (.A(_06138_),
    .B(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__a32o_1 _11097_ (.A1(\cur_mb_mem[165][7] ),
    .A2(_06137_),
    .A3(_06132_),
    .B1(_06141_),
    .B2(\cur_mb_mem[118][7] ),
    .X(_06142_));
 sky130_fd_sc_hd__buf_4 _11098_ (.A(_06022_),
    .X(_06143_));
 sky130_fd_sc_hd__and2_4 _11099_ (.A(_06140_),
    .B(_06143_),
    .X(_06144_));
 sky130_fd_sc_hd__a32o_2 _11100_ (.A1(\cur_mb_mem[148][7] ),
    .A2(_06134_),
    .A3(_05978_),
    .B1(_06144_),
    .B2(\cur_mb_mem[70][7] ),
    .X(_06145_));
 sky130_fd_sc_hd__buf_12 _11101_ (.A(net246),
    .X(_06146_));
 sky130_fd_sc_hd__clkbuf_16 _11102_ (.A(_06130_),
    .X(_06147_));
 sky130_fd_sc_hd__and2_4 _11103_ (.A(_06146_),
    .B(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__clkbuf_8 _11104_ (.A(_06099_),
    .X(_06149_));
 sky130_fd_sc_hd__buf_6 _11105_ (.A(_05940_),
    .X(_06150_));
 sky130_fd_sc_hd__and2_4 _11106_ (.A(_06149_),
    .B(_06150_),
    .X(_06151_));
 sky130_fd_sc_hd__clkbuf_8 _11107_ (.A(_05977_),
    .X(_06152_));
 sky130_fd_sc_hd__buf_8 _11108_ (.A(_06130_),
    .X(_06153_));
 sky130_fd_sc_hd__and3_2 _11109_ (.A(\cur_mb_mem[149][7] ),
    .B(_06152_),
    .C(_06153_),
    .X(_06154_));
 sky130_fd_sc_hd__a221o_1 _11110_ (.A1(\cur_mb_mem[133][7] ),
    .A2(_06148_),
    .B1(_06151_),
    .B2(\cur_mb_mem[223][7] ),
    .C1(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__or3_1 _11111_ (.A(_06142_),
    .B(_06145_),
    .C(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__and2_2 _11112_ (.A(_06112_),
    .B(_06132_),
    .X(_06157_));
 sky130_fd_sc_hd__clkbuf_8 _11113_ (.A(_04429_),
    .X(_06158_));
 sky130_fd_sc_hd__buf_12 _11114_ (.A(_06139_),
    .X(_06159_));
 sky130_fd_sc_hd__and2_4 _11115_ (.A(_06158_),
    .B(_06159_),
    .X(_06160_));
 sky130_fd_sc_hd__or4b_4 _11116_ (.A(_04653_),
    .B(_04458_),
    .C(_04692_),
    .D_N(_04669_),
    .X(_06161_));
 sky130_fd_sc_hd__nor2_8 _11117_ (.A(_06161_),
    .B(_05899_),
    .Y(_06162_));
 sky130_fd_sc_hd__a32o_2 _11118_ (.A1(\cur_mb_mem[20][7] ),
    .A2(_06134_),
    .A3(_05975_),
    .B1(_06162_),
    .B2(\cur_mb_mem[4][7] ),
    .X(_06163_));
 sky130_fd_sc_hd__a221o_1 _11119_ (.A1(\cur_mb_mem[5][7] ),
    .A2(_06157_),
    .B1(_06160_),
    .B2(\cur_mb_mem[246][7] ),
    .C1(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__buf_6 _11120_ (.A(_04429_),
    .X(_06165_));
 sky130_fd_sc_hd__buf_12 _11121_ (.A(net265),
    .X(_06166_));
 sky130_fd_sc_hd__and2_4 _11122_ (.A(_06165_),
    .B(_06166_),
    .X(_06167_));
 sky130_fd_sc_hd__a32o_2 _11123_ (.A1(\cur_mb_mem[213][7] ),
    .A2(_05942_),
    .A3(_06133_),
    .B1(_06167_),
    .B2(\cur_mb_mem[244][7] ),
    .X(_06168_));
 sky130_fd_sc_hd__or4_2 _11124_ (.A(_06136_),
    .B(_06156_),
    .C(_06164_),
    .D(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__clkbuf_8 _11125_ (.A(_05055_),
    .X(_06170_));
 sky130_fd_sc_hd__clkbuf_16 _11126_ (.A(net223),
    .X(_06171_));
 sky130_fd_sc_hd__and2_4 _11127_ (.A(_06170_),
    .B(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__a32o_1 _11128_ (.A1(\cur_mb_mem[63][7] ),
    .A2(_04424_),
    .A3(_05058_),
    .B1(_06172_),
    .B2(\cur_mb_mem[50][7] ),
    .X(_06173_));
 sky130_fd_sc_hd__and2_4 _11129_ (.A(_06099_),
    .B(_05977_),
    .X(_06174_));
 sky130_fd_sc_hd__a32o_1 _11130_ (.A1(\cur_mb_mem[207][7] ),
    .A2(_04424_),
    .A3(_06094_),
    .B1(_06174_),
    .B2(\cur_mb_mem[159][7] ),
    .X(_06175_));
 sky130_fd_sc_hd__nand4_4 _11131_ (.A(_04654_),
    .B(_04459_),
    .C(_04670_),
    .D(_04692_),
    .Y(_06176_));
 sky130_fd_sc_hd__or4b_4 _11132_ (.A(_04426_),
    .B(_04427_),
    .C(_04428_),
    .D_N(_04425_),
    .X(_06177_));
 sky130_fd_sc_hd__nor2_8 _11133_ (.A(net221),
    .B(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__clkbuf_16 _11134_ (.A(_06095_),
    .X(_06179_));
 sky130_fd_sc_hd__and2_4 _11135_ (.A(_06179_),
    .B(_05997_),
    .X(_06180_));
 sky130_fd_sc_hd__and3_1 _11136_ (.A(\cur_mb_mem[160][7] ),
    .B(_05923_),
    .C(_05971_),
    .X(_06181_));
 sky130_fd_sc_hd__a31o_1 _11137_ (.A1(\cur_mb_mem[64][7] ),
    .A2(_06024_),
    .A3(_05972_),
    .B1(_06181_),
    .X(_06182_));
 sky130_fd_sc_hd__a221o_1 _11138_ (.A1(\cur_mb_mem[31][7] ),
    .A2(_06178_),
    .B1(_06180_),
    .B2(\cur_mb_mem[231][7] ),
    .C1(_06182_),
    .X(_06183_));
 sky130_fd_sc_hd__or4_1 _11139_ (.A(_06169_),
    .B(_06173_),
    .C(_06175_),
    .D(_06183_),
    .X(_06184_));
 sky130_fd_sc_hd__nor2_8 _11140_ (.A(_05897_),
    .B(_05906_),
    .Y(_06185_));
 sky130_fd_sc_hd__buf_6 _11141_ (.A(_06139_),
    .X(_06186_));
 sky130_fd_sc_hd__buf_8 _11142_ (.A(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__buf_4 _11143_ (.A(_05977_),
    .X(_06188_));
 sky130_fd_sc_hd__and2_4 _11144_ (.A(_06159_),
    .B(_06188_),
    .X(_06189_));
 sky130_fd_sc_hd__a32o_1 _11145_ (.A1(\cur_mb_mem[214][7] ),
    .A2(_06187_),
    .A3(_05942_),
    .B1(_06189_),
    .B2(\cur_mb_mem[150][7] ),
    .X(_06190_));
 sky130_fd_sc_hd__buf_12 _11146_ (.A(_06159_),
    .X(_06191_));
 sky130_fd_sc_hd__buf_8 _11147_ (.A(_05921_),
    .X(_06192_));
 sky130_fd_sc_hd__and2_4 _11148_ (.A(_06191_),
    .B(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__a32o_1 _11149_ (.A1(\cur_mb_mem[86][7] ),
    .A2(_05925_),
    .A3(_06187_),
    .B1(_06193_),
    .B2(\cur_mb_mem[166][7] ),
    .X(_06194_));
 sky130_fd_sc_hd__and2_4 _11150_ (.A(_06026_),
    .B(_05921_),
    .X(_06195_));
 sky130_fd_sc_hd__nor2_8 _11151_ (.A(_06161_),
    .B(_05965_),
    .Y(_06196_));
 sky130_fd_sc_hd__a22o_2 _11152_ (.A1(\cur_mb_mem[164][7] ),
    .A2(_06195_),
    .B1(net220),
    .B2(\cur_mb_mem[132][7] ),
    .X(_06197_));
 sky130_fd_sc_hd__clkbuf_8 _11153_ (.A(_05055_),
    .X(_06198_));
 sky130_fd_sc_hd__clkbuf_16 _11154_ (.A(_06139_),
    .X(_06199_));
 sky130_fd_sc_hd__and3_1 _11155_ (.A(\cur_mb_mem[54][7] ),
    .B(_06198_),
    .C(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__a31o_1 _11156_ (.A1(\cur_mb_mem[196][7] ),
    .A2(_05890_),
    .A3(_06091_),
    .B1(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__buf_12 _11157_ (.A(_05926_),
    .X(_06202_));
 sky130_fd_sc_hd__and2_4 _11158_ (.A(_06202_),
    .B(_06140_),
    .X(_06203_));
 sky130_fd_sc_hd__buf_12 _11159_ (.A(_06159_),
    .X(_06204_));
 sky130_fd_sc_hd__and2_4 _11160_ (.A(_06204_),
    .B(_06019_),
    .X(_06205_));
 sky130_fd_sc_hd__a22o_1 _11161_ (.A1(\cur_mb_mem[6][7] ),
    .A2(_06203_),
    .B1(_06205_),
    .B2(\cur_mb_mem[182][7] ),
    .X(_06206_));
 sky130_fd_sc_hd__clkbuf_8 _11162_ (.A(_06050_),
    .X(_06207_));
 sky130_fd_sc_hd__buf_8 _11163_ (.A(_06130_),
    .X(_06208_));
 sky130_fd_sc_hd__and2_4 _11164_ (.A(_06207_),
    .B(_06208_),
    .X(_06209_));
 sky130_fd_sc_hd__buf_12 _11165_ (.A(_06139_),
    .X(_06210_));
 sky130_fd_sc_hd__and2_4 _11166_ (.A(_06210_),
    .B(_05933_),
    .X(_06211_));
 sky130_fd_sc_hd__a22o_1 _11167_ (.A1(\cur_mb_mem[117][7] ),
    .A2(_06209_),
    .B1(_06211_),
    .B2(\cur_mb_mem[134][7] ),
    .X(_06212_));
 sky130_fd_sc_hd__or4_1 _11168_ (.A(_06197_),
    .B(_06201_),
    .C(_06206_),
    .D(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__or4_1 _11169_ (.A(_06185_),
    .B(_06190_),
    .C(_06194_),
    .D(_06213_),
    .X(_06214_));
 sky130_fd_sc_hd__buf_12 _11170_ (.A(net263),
    .X(_06215_));
 sky130_fd_sc_hd__buf_12 _11171_ (.A(_06018_),
    .X(_06216_));
 sky130_fd_sc_hd__and2_4 _11172_ (.A(_06215_),
    .B(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__and2_4 _11173_ (.A(_06023_),
    .B(_06132_),
    .X(_06218_));
 sky130_fd_sc_hd__a22o_4 _11174_ (.A1(\cur_mb_mem[180][7] ),
    .A2(_06217_),
    .B1(_06218_),
    .B2(\cur_mb_mem[69][7] ),
    .X(_06219_));
 sky130_fd_sc_hd__buf_12 _11175_ (.A(_06130_),
    .X(_06220_));
 sky130_fd_sc_hd__and2_4 _11176_ (.A(_06170_),
    .B(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__a32o_1 _11177_ (.A1(\cur_mb_mem[181][7] ),
    .A2(_06037_),
    .A3(_06133_),
    .B1(_06221_),
    .B2(\cur_mb_mem[53][7] ),
    .X(_06222_));
 sky130_fd_sc_hd__buf_12 _11178_ (.A(_06134_),
    .X(_06223_));
 sky130_fd_sc_hd__buf_4 _11179_ (.A(_05997_),
    .X(_06224_));
 sky130_fd_sc_hd__and3_1 _11180_ (.A(\cur_mb_mem[229][7] ),
    .B(_06132_),
    .C(_06224_),
    .X(_06225_));
 sky130_fd_sc_hd__a31o_1 _11181_ (.A1(\cur_mb_mem[228][7] ),
    .A2(_06223_),
    .A3(_06066_),
    .B1(_06225_),
    .X(_06226_));
 sky130_fd_sc_hd__and3_1 _11182_ (.A(\cur_mb_mem[230][7] ),
    .B(_06186_),
    .C(_06224_),
    .X(_06227_));
 sky130_fd_sc_hd__a31o_1 _11183_ (.A1(\cur_mb_mem[245][7] ),
    .A2(_04431_),
    .A3(_06133_),
    .B1(_06227_),
    .X(_06228_));
 sky130_fd_sc_hd__or4_4 _11184_ (.A(_06219_),
    .B(_06222_),
    .C(_06226_),
    .D(_06228_),
    .X(_06229_));
 sky130_fd_sc_hd__buf_8 _11185_ (.A(net253),
    .X(_06230_));
 sky130_fd_sc_hd__and2_4 _11186_ (.A(_06230_),
    .B(_06147_),
    .X(_06231_));
 sky130_fd_sc_hd__buf_8 _11187_ (.A(net2008),
    .X(_06232_));
 sky130_fd_sc_hd__buf_4 _11188_ (.A(_06022_),
    .X(_06233_));
 sky130_fd_sc_hd__and2_4 _11189_ (.A(_06232_),
    .B(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__clkbuf_16 _11190_ (.A(net233),
    .X(_06235_));
 sky130_fd_sc_hd__and2_4 _11191_ (.A(_06235_),
    .B(_06147_),
    .X(_06236_));
 sky130_fd_sc_hd__a32o_1 _11192_ (.A1(\cur_mb_mem[198][7] ),
    .A2(_06187_),
    .A3(_06093_),
    .B1(_06236_),
    .B2(\cur_mb_mem[21][7] ),
    .X(_06237_));
 sky130_fd_sc_hd__a221o_1 _11193_ (.A1(\cur_mb_mem[85][7] ),
    .A2(_06231_),
    .B1(_06234_),
    .B2(\cur_mb_mem[68][7] ),
    .C1(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__and2_4 _11194_ (.A(_05890_),
    .B(_06052_),
    .X(_06239_));
 sky130_fd_sc_hd__buf_6 _11195_ (.A(_05055_),
    .X(_06240_));
 sky130_fd_sc_hd__and2_4 _11196_ (.A(_06240_),
    .B(_06232_),
    .X(_06241_));
 sky130_fd_sc_hd__and2_4 _11197_ (.A(_06204_),
    .B(_06235_),
    .X(_06242_));
 sky130_fd_sc_hd__a32o_1 _11198_ (.A1(\cur_mb_mem[84][7] ),
    .A2(_06223_),
    .A3(_05925_),
    .B1(_06242_),
    .B2(\cur_mb_mem[22][7] ),
    .X(_06243_));
 sky130_fd_sc_hd__a221o_2 _11199_ (.A1(\cur_mb_mem[116][7] ),
    .A2(_06239_),
    .B1(_06241_),
    .B2(\cur_mb_mem[52][7] ),
    .C1(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__or4_1 _11200_ (.A(_06214_),
    .B(_06229_),
    .C(_06238_),
    .D(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__clkbuf_8 _11201_ (.A(_05944_),
    .X(_06246_));
 sky130_fd_sc_hd__clkbuf_4 _11202_ (.A(_05997_),
    .X(_06247_));
 sky130_fd_sc_hd__and2_4 _11203_ (.A(_06246_),
    .B(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__a32o_1 _11204_ (.A1(\cur_mb_mem[167][7] ),
    .A2(_05923_),
    .A3(_06097_),
    .B1(_06248_),
    .B2(\cur_mb_mem[237][7] ),
    .X(_06249_));
 sky130_fd_sc_hd__and2_4 _11205_ (.A(_06033_),
    .B(_05933_),
    .X(_06250_));
 sky130_fd_sc_hd__buf_12 _11206_ (.A(net228),
    .X(_06251_));
 sky130_fd_sc_hd__and2_4 _11207_ (.A(_06152_),
    .B(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__a22o_2 _11208_ (.A1(\cur_mb_mem[141][7] ),
    .A2(_06250_),
    .B1(_06252_),
    .B2(\cur_mb_mem[145][7] ),
    .X(_06253_));
 sky130_fd_sc_hd__clkbuf_16 _11209_ (.A(net222),
    .X(_06254_));
 sky130_fd_sc_hd__clkbuf_4 _11210_ (.A(_05997_),
    .X(_06255_));
 sky130_fd_sc_hd__and2_4 _11211_ (.A(_06254_),
    .B(_06255_),
    .X(_06256_));
 sky130_fd_sc_hd__or4b_1 _11212_ (.A(_04425_),
    .B(_04427_),
    .C(_04428_),
    .D_N(_04426_),
    .X(_06257_));
 sky130_fd_sc_hd__buf_8 _11213_ (.A(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__nor2_8 _11214_ (.A(net221),
    .B(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__a22o_1 _11215_ (.A1(\cur_mb_mem[226][7] ),
    .A2(_06256_),
    .B1(_06259_),
    .B2(\cur_mb_mem[47][7] ),
    .X(_06260_));
 sky130_fd_sc_hd__buf_8 _11216_ (.A(_05917_),
    .X(_06261_));
 sky130_fd_sc_hd__and3_1 _11217_ (.A(\cur_mb_mem[235][7] ),
    .B(_06261_),
    .C(_06066_),
    .X(_06262_));
 sky130_fd_sc_hd__a31o_1 _11218_ (.A1(\cur_mb_mem[247][7] ),
    .A2(_04431_),
    .A3(_06098_),
    .B1(_06262_),
    .X(_06263_));
 sky130_fd_sc_hd__or4_1 _11219_ (.A(_06249_),
    .B(_06253_),
    .C(_06260_),
    .D(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__or4b_4 _11220_ (.A(_04459_),
    .B(_04670_),
    .C(_04692_),
    .D_N(_04654_),
    .X(_06265_));
 sky130_fd_sc_hd__nor2_2 _11221_ (.A(_06265_),
    .B(_05965_),
    .Y(_06266_));
 sky130_fd_sc_hd__buf_4 _11222_ (.A(_05983_),
    .X(_06267_));
 sky130_fd_sc_hd__clkbuf_8 _11223_ (.A(_06267_),
    .X(_06268_));
 sky130_fd_sc_hd__and2_4 _11224_ (.A(_06268_),
    .B(_06208_),
    .X(_06269_));
 sky130_fd_sc_hd__clkbuf_8 _11225_ (.A(_05940_),
    .X(_06270_));
 sky130_fd_sc_hd__and2_4 _11226_ (.A(_06270_),
    .B(_05995_),
    .X(_06271_));
 sky130_fd_sc_hd__a32o_4 _11227_ (.A1(\cur_mb_mem[252][7] ),
    .A2(_04431_),
    .A3(_05938_),
    .B1(_06271_),
    .B2(\cur_mb_mem[209][7] ),
    .X(_06272_));
 sky130_fd_sc_hd__a221o_1 _11228_ (.A1(\cur_mb_mem[130][7] ),
    .A2(_06266_),
    .B1(_06269_),
    .B2(\cur_mb_mem[101][7] ),
    .C1(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__and3_1 _11229_ (.A(\cur_mb_mem[13][7] ),
    .B(_06113_),
    .C(_05961_),
    .X(_06274_));
 sky130_fd_sc_hd__a31o_1 _11230_ (.A1(\cur_mb_mem[62][7] ),
    .A2(_05059_),
    .A3(_06025_),
    .B1(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__or4b_4 _11231_ (.A(_04653_),
    .B(_04458_),
    .C(_04670_),
    .D_N(_04692_),
    .X(_06276_));
 sky130_fd_sc_hd__nor2_4 _11232_ (.A(_05899_),
    .B(_06276_),
    .Y(_06277_));
 sky130_fd_sc_hd__a32o_1 _11233_ (.A1(\cur_mb_mem[206][7] ),
    .A2(_06025_),
    .A3(_06094_),
    .B1(_06277_),
    .B2(\cur_mb_mem[8][7] ),
    .X(_06278_));
 sky130_fd_sc_hd__or4_1 _11234_ (.A(_06264_),
    .B(_06273_),
    .C(_06275_),
    .D(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__and2_4 _11235_ (.A(_06254_),
    .B(_06138_),
    .X(_06280_));
 sky130_fd_sc_hd__and2_1 _11236_ (.A(_06060_),
    .B(_05974_),
    .X(_06281_));
 sky130_fd_sc_hd__clkbuf_16 _11237_ (.A(_06281_),
    .X(_06282_));
 sky130_fd_sc_hd__clkbuf_8 _11238_ (.A(_06079_),
    .X(_06283_));
 sky130_fd_sc_hd__and2_4 _11239_ (.A(_06283_),
    .B(_05922_),
    .X(_06284_));
 sky130_fd_sc_hd__nor2_8 _11240_ (.A(_06276_),
    .B(_06177_),
    .Y(_06285_));
 sky130_fd_sc_hd__a22o_1 _11241_ (.A1(\cur_mb_mem[162][7] ),
    .A2(_06284_),
    .B1(_06285_),
    .B2(\cur_mb_mem[24][7] ),
    .X(_06286_));
 sky130_fd_sc_hd__a221o_1 _11242_ (.A1(\cur_mb_mem[114][7] ),
    .A2(_06280_),
    .B1(_06282_),
    .B2(\cur_mb_mem[19][7] ),
    .C1(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__and2_4 _11243_ (.A(_05895_),
    .B(_06022_),
    .X(_06288_));
 sky130_fd_sc_hd__buf_8 _11244_ (.A(_06060_),
    .X(_06289_));
 sky130_fd_sc_hd__and2_4 _11245_ (.A(_06202_),
    .B(_06289_),
    .X(_06290_));
 sky130_fd_sc_hd__nor2_4 _11246_ (.A(_06258_),
    .B(_05963_),
    .Y(_06291_));
 sky130_fd_sc_hd__nor2_8 _11247_ (.A(_06276_),
    .B(_05965_),
    .Y(_06292_));
 sky130_fd_sc_hd__a22o_1 _11248_ (.A1(\cur_mb_mem[33][7] ),
    .A2(_06291_),
    .B1(_06292_),
    .B2(\cur_mb_mem[136][7] ),
    .X(_06293_));
 sky130_fd_sc_hd__a221o_2 _11249_ (.A1(\cur_mb_mem[72][7] ),
    .A2(_06288_),
    .B1(_06290_),
    .B2(\cur_mb_mem[3][7] ),
    .C1(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__nor2_8 _11250_ (.A(_06176_),
    .B(_05899_),
    .Y(_06295_));
 sky130_fd_sc_hd__nand2_4 _11251_ (.A(_04969_),
    .B(_05112_),
    .Y(_06296_));
 sky130_fd_sc_hd__nor2_4 _11252_ (.A(net221),
    .B(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__buf_8 _11253_ (.A(_06267_),
    .X(_06298_));
 sky130_fd_sc_hd__buf_8 _11254_ (.A(_06298_),
    .X(_06299_));
 sky130_fd_sc_hd__buf_8 _11255_ (.A(net252),
    .X(_06300_));
 sky130_fd_sc_hd__and2_4 _11256_ (.A(_06300_),
    .B(_06003_),
    .X(_06301_));
 sky130_fd_sc_hd__a32o_1 _11257_ (.A1(\cur_mb_mem[96][7] ),
    .A2(_06299_),
    .A3(_05972_),
    .B1(_06301_),
    .B2(\cur_mb_mem[11][7] ),
    .X(_06302_));
 sky130_fd_sc_hd__a221o_1 _11258_ (.A1(\cur_mb_mem[15][7] ),
    .A2(_06295_),
    .B1(_06297_),
    .B2(\cur_mb_mem[95][7] ),
    .C1(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__and2_4 _11259_ (.A(_06068_),
    .B(_06032_),
    .X(_06304_));
 sky130_fd_sc_hd__nor2_8 _11260_ (.A(net221),
    .B(_05965_),
    .Y(_06305_));
 sky130_fd_sc_hd__and3_1 _11261_ (.A(\cur_mb_mem[103][7] ),
    .B(_06298_),
    .C(_06097_),
    .X(_06306_));
 sky130_fd_sc_hd__a31o_1 _11262_ (.A1(\cur_mb_mem[55][7] ),
    .A2(_05058_),
    .A3(_06098_),
    .B1(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__a221o_1 _11263_ (.A1(\cur_mb_mem[255][7] ),
    .A2(_06304_),
    .B1(_06305_),
    .B2(\cur_mb_mem[143][7] ),
    .C1(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__or4_1 _11264_ (.A(_06287_),
    .B(_06294_),
    .C(_06303_),
    .D(_06308_),
    .X(_06309_));
 sky130_fd_sc_hd__or4_1 _11265_ (.A(_06184_),
    .B(_06245_),
    .C(_06279_),
    .D(_06309_),
    .X(_06310_));
 sky130_fd_sc_hd__or4_4 _11266_ (.A(_06043_),
    .B(_06090_),
    .C(_06129_),
    .D(_06310_),
    .X(_06311_));
 sky130_fd_sc_hd__clkbuf_16 _11267_ (.A(_05917_),
    .X(_06312_));
 sky130_fd_sc_hd__buf_4 _11268_ (.A(_05983_),
    .X(_06313_));
 sky130_fd_sc_hd__and2_2 _11269_ (.A(_06312_),
    .B(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__buf_8 _11270_ (.A(net236),
    .X(_06315_));
 sky130_fd_sc_hd__and2_4 _11271_ (.A(_06036_),
    .B(_06315_),
    .X(_06316_));
 sky130_fd_sc_hd__and2_4 _11272_ (.A(_05896_),
    .B(_05941_),
    .X(_06317_));
 sky130_fd_sc_hd__nor2_8 _11273_ (.A(_05963_),
    .B(_06177_),
    .Y(_06318_));
 sky130_fd_sc_hd__a22o_1 _11274_ (.A1(\cur_mb_mem[216][7] ),
    .A2(_06317_),
    .B1(_06318_),
    .B2(\cur_mb_mem[17][7] ),
    .X(_06319_));
 sky130_fd_sc_hd__a221o_1 _11275_ (.A1(\cur_mb_mem[107][7] ),
    .A2(_06314_),
    .B1(_06316_),
    .B2(\cur_mb_mem[176][7] ),
    .C1(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__buf_8 _11276_ (.A(_05900_),
    .X(_06321_));
 sky130_fd_sc_hd__and2_4 _11277_ (.A(_06321_),
    .B(_06027_),
    .X(_06322_));
 sky130_fd_sc_hd__a32o_1 _11278_ (.A1(\cur_mb_mem[243][7] ),
    .A2(_04432_),
    .A3(_06064_),
    .B1(_06322_),
    .B2(\cur_mb_mem[108][7] ),
    .X(_06323_));
 sky130_fd_sc_hd__buf_4 _11279_ (.A(_06081_),
    .X(_06324_));
 sky130_fd_sc_hd__and2_4 _11280_ (.A(_06312_),
    .B(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__a32o_1 _11281_ (.A1(\cur_mb_mem[208][7] ),
    .A2(_06106_),
    .A3(_05973_),
    .B1(_06325_),
    .B2(\cur_mb_mem[203][7] ),
    .X(_06326_));
 sky130_fd_sc_hd__clkbuf_16 _11282_ (.A(_05892_),
    .X(_06327_));
 sky130_fd_sc_hd__and2_4 _11283_ (.A(_06327_),
    .B(_06121_),
    .X(_06328_));
 sky130_fd_sc_hd__a32o_2 _11284_ (.A1(\cur_mb_mem[75][7] ),
    .A2(_06049_),
    .A3(_06024_),
    .B1(_06328_),
    .B2(\cur_mb_mem[73][7] ),
    .X(_06329_));
 sky130_fd_sc_hd__and2_4 _11285_ (.A(_06171_),
    .B(_06027_),
    .X(_06330_));
 sky130_fd_sc_hd__a32o_1 _11286_ (.A1(\cur_mb_mem[218][7] ),
    .A2(_06035_),
    .A3(_06106_),
    .B1(_06330_),
    .B2(\cur_mb_mem[98][7] ),
    .X(_06331_));
 sky130_fd_sc_hd__or4_4 _11287_ (.A(_06323_),
    .B(_06326_),
    .C(_06329_),
    .D(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__clkbuf_8 _11288_ (.A(_05920_),
    .X(_06333_));
 sky130_fd_sc_hd__and2_4 _11289_ (.A(_06076_),
    .B(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__and2_4 _11290_ (.A(_04430_),
    .B(_06283_),
    .X(_06335_));
 sky130_fd_sc_hd__clkbuf_8 _11291_ (.A(_05911_),
    .X(_06336_));
 sky130_fd_sc_hd__and3_1 _11292_ (.A(\cur_mb_mem[188][7] ),
    .B(_05937_),
    .C(_06036_),
    .X(_06337_));
 sky130_fd_sc_hd__a31o_1 _11293_ (.A1(\cur_mb_mem[217][7] ),
    .A2(_06336_),
    .A3(_05942_),
    .B1(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__a221o_1 _11294_ (.A1(\cur_mb_mem[161][7] ),
    .A2(_06334_),
    .B1(_06335_),
    .B2(\cur_mb_mem[242][7] ),
    .C1(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__and2_2 _11295_ (.A(_05902_),
    .B(_06057_),
    .X(_06340_));
 sky130_fd_sc_hd__buf_12 _11296_ (.A(net222),
    .X(_06341_));
 sky130_fd_sc_hd__and2_4 _11297_ (.A(_06341_),
    .B(_06270_),
    .X(_06342_));
 sky130_fd_sc_hd__buf_8 _11298_ (.A(net226),
    .X(_06343_));
 sky130_fd_sc_hd__and2_4 _11299_ (.A(_06343_),
    .B(_06147_),
    .X(_06344_));
 sky130_fd_sc_hd__a32o_1 _11300_ (.A1(\cur_mb_mem[241][7] ),
    .A2(_04431_),
    .A3(_05994_),
    .B1(_06344_),
    .B2(\cur_mb_mem[37][7] ),
    .X(_06345_));
 sky130_fd_sc_hd__a221o_1 _11301_ (.A1(\cur_mb_mem[76][7] ),
    .A2(_06340_),
    .B1(_06342_),
    .B2(\cur_mb_mem[210][7] ),
    .C1(_06345_),
    .X(_06346_));
 sky130_fd_sc_hd__buf_12 _11302_ (.A(_06060_),
    .X(_06347_));
 sky130_fd_sc_hd__buf_4 _11303_ (.A(_05939_),
    .X(_06348_));
 sky130_fd_sc_hd__and2_4 _11304_ (.A(_06347_),
    .B(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__clkbuf_8 _11305_ (.A(_05055_),
    .X(_06350_));
 sky130_fd_sc_hd__and2_4 _11306_ (.A(_06350_),
    .B(_05895_),
    .X(_06351_));
 sky130_fd_sc_hd__buf_4 _11307_ (.A(_06081_),
    .X(_06352_));
 sky130_fd_sc_hd__buf_12 _11308_ (.A(net227),
    .X(_06353_));
 sky130_fd_sc_hd__and2_4 _11309_ (.A(_06352_),
    .B(_06353_),
    .X(_06354_));
 sky130_fd_sc_hd__buf_12 _11310_ (.A(_06060_),
    .X(_06355_));
 sky130_fd_sc_hd__and2_2 _11311_ (.A(_06355_),
    .B(_06039_),
    .X(_06356_));
 sky130_fd_sc_hd__a22o_1 _11312_ (.A1(\cur_mb_mem[193][7] ),
    .A2(_06354_),
    .B1(_06356_),
    .B2(\cur_mb_mem[179][7] ),
    .X(_06357_));
 sky130_fd_sc_hd__a221o_1 _11313_ (.A1(\cur_mb_mem[211][7] ),
    .A2(_06349_),
    .B1(_06351_),
    .B2(\cur_mb_mem[56][7] ),
    .C1(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__and2_4 _11314_ (.A(_06170_),
    .B(_06011_),
    .X(_06359_));
 sky130_fd_sc_hd__nor2_8 _11315_ (.A(_06161_),
    .B(_06258_),
    .Y(_06360_));
 sky130_fd_sc_hd__and2_4 _11316_ (.A(_06003_),
    .B(_06008_),
    .X(_06361_));
 sky130_fd_sc_hd__a32o_1 _11317_ (.A1(\cur_mb_mem[59][7] ),
    .A2(_05058_),
    .A3(_06049_),
    .B1(_06361_),
    .B2(\cur_mb_mem[91][7] ),
    .X(_06362_));
 sky130_fd_sc_hd__a221o_1 _11318_ (.A1(\cur_mb_mem[61][7] ),
    .A2(_06359_),
    .B1(_06360_),
    .B2(\cur_mb_mem[36][7] ),
    .C1(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__or4_1 _11319_ (.A(_06339_),
    .B(_06346_),
    .C(_06358_),
    .D(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__clkbuf_16 _11320_ (.A(_05926_),
    .X(_06365_));
 sky130_fd_sc_hd__buf_8 _11321_ (.A(_05952_),
    .X(_06366_));
 sky130_fd_sc_hd__and2_4 _11322_ (.A(_06365_),
    .B(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__and2_4 _11323_ (.A(_06171_),
    .B(_06143_),
    .X(_06368_));
 sky130_fd_sc_hd__a22o_1 _11324_ (.A1(\cur_mb_mem[14][7] ),
    .A2(_06367_),
    .B1(_06368_),
    .B2(\cur_mb_mem[66][7] ),
    .X(_06369_));
 sky130_fd_sc_hd__and2_1 _11325_ (.A(_06246_),
    .B(_06091_),
    .X(_06370_));
 sky130_fd_sc_hd__a32o_2 _11326_ (.A1(\cur_mb_mem[254][7] ),
    .A2(_04432_),
    .A3(_06025_),
    .B1(_06370_),
    .B2(\cur_mb_mem[205][7] ),
    .X(_06371_));
 sky130_fd_sc_hd__clkbuf_16 _11327_ (.A(_06095_),
    .X(_06372_));
 sky130_fd_sc_hd__and2_4 _11328_ (.A(_06343_),
    .B(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__a32o_1 _11329_ (.A1(\cur_mb_mem[147][7] ),
    .A2(_06064_),
    .A3(_05980_),
    .B1(_06373_),
    .B2(\cur_mb_mem[39][7] ),
    .X(_06374_));
 sky130_fd_sc_hd__and3_1 _11330_ (.A(\cur_mb_mem[2][7] ),
    .B(_06113_),
    .C(_06283_),
    .X(_06375_));
 sky130_fd_sc_hd__a31o_1 _11331_ (.A1(\cur_mb_mem[51][7] ),
    .A2(_05059_),
    .A3(_06064_),
    .B1(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__or4_1 _11332_ (.A(_06369_),
    .B(_06371_),
    .C(_06374_),
    .D(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__buf_4 _11333_ (.A(net253),
    .X(_06378_));
 sky130_fd_sc_hd__and2_4 _11334_ (.A(_06378_),
    .B(_06355_),
    .X(_06379_));
 sky130_fd_sc_hd__buf_12 _11335_ (.A(_06079_),
    .X(_06380_));
 sky130_fd_sc_hd__and2_4 _11336_ (.A(_06380_),
    .B(_06152_),
    .X(_06381_));
 sky130_fd_sc_hd__buf_8 _11337_ (.A(net249),
    .X(_06382_));
 sky130_fd_sc_hd__and2_4 _11338_ (.A(_06289_),
    .B(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__a32o_2 _11339_ (.A1(\cur_mb_mem[163][7] ),
    .A2(_06064_),
    .A3(_05956_),
    .B1(_06383_),
    .B2(\cur_mb_mem[131][7] ),
    .X(_06384_));
 sky130_fd_sc_hd__a221o_1 _11340_ (.A1(\cur_mb_mem[83][7] ),
    .A2(_06379_),
    .B1(_06381_),
    .B2(\cur_mb_mem[146][7] ),
    .C1(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__and2_2 _11341_ (.A(_06283_),
    .B(_06037_),
    .X(_06386_));
 sky130_fd_sc_hd__buf_8 _11342_ (.A(_05917_),
    .X(_06387_));
 sky130_fd_sc_hd__and2_4 _11343_ (.A(_06387_),
    .B(_06146_),
    .X(_06388_));
 sky130_fd_sc_hd__and3_1 _11344_ (.A(\cur_mb_mem[82][7] ),
    .B(_06283_),
    .C(_05916_),
    .X(_06389_));
 sky130_fd_sc_hd__a31o_1 _11345_ (.A1(\cur_mb_mem[202][7] ),
    .A2(_06035_),
    .A3(_06094_),
    .B1(_06389_),
    .X(_06390_));
 sky130_fd_sc_hd__a221o_1 _11346_ (.A1(\cur_mb_mem[178][7] ),
    .A2(_06386_),
    .B1(_06388_),
    .B2(\cur_mb_mem[139][7] ),
    .C1(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__or4_1 _11347_ (.A(_06364_),
    .B(_06377_),
    .C(_06385_),
    .D(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__nor2_8 _11348_ (.A(_06265_),
    .B(_06258_),
    .Y(_06393_));
 sky130_fd_sc_hd__and2_4 _11349_ (.A(_05895_),
    .B(_06188_),
    .X(_06394_));
 sky130_fd_sc_hd__buf_8 _11350_ (.A(net225),
    .X(_06395_));
 sky130_fd_sc_hd__and2_4 _11351_ (.A(_06395_),
    .B(_06210_),
    .X(_06396_));
 sky130_fd_sc_hd__a32o_1 _11352_ (.A1(\cur_mb_mem[157][7] ),
    .A2(_05961_),
    .A3(_05980_),
    .B1(_06396_),
    .B2(\cur_mb_mem[38][7] ),
    .X(_06397_));
 sky130_fd_sc_hd__a221o_1 _11353_ (.A1(\cur_mb_mem[34][7] ),
    .A2(_06393_),
    .B1(_06394_),
    .B2(\cur_mb_mem[152][7] ),
    .C1(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__and2_4 _11354_ (.A(_06321_),
    .B(_06005_),
    .X(_06399_));
 sky130_fd_sc_hd__clkbuf_16 _11355_ (.A(_05917_),
    .X(_06400_));
 sky130_fd_sc_hd__clkbuf_8 _11356_ (.A(_05977_),
    .X(_06401_));
 sky130_fd_sc_hd__and2_4 _11357_ (.A(_06400_),
    .B(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__buf_4 _11358_ (.A(net232),
    .X(_06403_));
 sky130_fd_sc_hd__and2_4 _11359_ (.A(_06011_),
    .B(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__a32o_1 _11360_ (.A1(\cur_mb_mem[124][7] ),
    .A2(_05989_),
    .A3(_06119_),
    .B1(_06404_),
    .B2(\cur_mb_mem[29][7] ),
    .X(_06405_));
 sky130_fd_sc_hd__a221o_1 _11361_ (.A1(\cur_mb_mem[44][7] ),
    .A2(_06399_),
    .B1(_06402_),
    .B2(\cur_mb_mem[155][7] ),
    .C1(_06405_),
    .X(_06406_));
 sky130_fd_sc_hd__and2_1 _11362_ (.A(net250),
    .B(_05904_),
    .X(_06407_));
 sky130_fd_sc_hd__buf_8 _11363_ (.A(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__a32o_1 _11364_ (.A1(\cur_mb_mem[9][7] ),
    .A2(_06113_),
    .A3(_06336_),
    .B1(_06408_),
    .B2(\cur_mb_mem[10][7] ),
    .X(_06409_));
 sky130_fd_sc_hd__and2_1 _11365_ (.A(_04429_),
    .B(net256),
    .X(_06410_));
 sky130_fd_sc_hd__buf_6 _11366_ (.A(_06410_),
    .X(_06411_));
 sky130_fd_sc_hd__a32o_1 _11367_ (.A1(\cur_mb_mem[99][7] ),
    .A2(_06298_),
    .A3(_06063_),
    .B1(_06411_),
    .B2(\cur_mb_mem[248][7] ),
    .X(_06412_));
 sky130_fd_sc_hd__buf_8 _11368_ (.A(_05983_),
    .X(_06413_));
 sky130_fd_sc_hd__and2_1 _11369_ (.A(_06413_),
    .B(_06186_),
    .X(_06414_));
 sky130_fd_sc_hd__a32o_1 _11370_ (.A1(\cur_mb_mem[105][7] ),
    .A2(_06336_),
    .A3(_06298_),
    .B1(_06414_),
    .B2(\cur_mb_mem[102][7] ),
    .X(_06415_));
 sky130_fd_sc_hd__and2_1 _11371_ (.A(_05904_),
    .B(net224),
    .X(_06416_));
 sky130_fd_sc_hd__buf_8 _11372_ (.A(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__a32o_1 _11373_ (.A1(\cur_mb_mem[121][7] ),
    .A2(_06336_),
    .A3(_06053_),
    .B1(_06417_),
    .B2(\cur_mb_mem[74][7] ),
    .X(_06418_));
 sky130_fd_sc_hd__or4_1 _11374_ (.A(_06409_),
    .B(_06412_),
    .C(_06415_),
    .D(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__or3_1 _11375_ (.A(_06398_),
    .B(_06406_),
    .C(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__and3_1 _11376_ (.A(\cur_mb_mem[125][7] ),
    .B(_05961_),
    .C(_06053_),
    .X(_06421_));
 sky130_fd_sc_hd__buf_12 _11377_ (.A(_05900_),
    .X(_06422_));
 sky130_fd_sc_hd__and2_4 _11378_ (.A(_06422_),
    .B(_05933_),
    .X(_06423_));
 sky130_fd_sc_hd__a32o_2 _11379_ (.A1(\cur_mb_mem[18][7] ),
    .A2(_06283_),
    .A3(_05976_),
    .B1(_06423_),
    .B2(\cur_mb_mem[140][7] ),
    .X(_06424_));
 sky130_fd_sc_hd__a311o_1 _11380_ (.A1(\cur_mb_mem[123][7] ),
    .A2(_06049_),
    .A3(_06119_),
    .B1(_06421_),
    .C1(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__buf_8 _11381_ (.A(_06137_),
    .X(_06426_));
 sky130_fd_sc_hd__and3_1 _11382_ (.A(\cur_mb_mem[170][7] ),
    .B(_05959_),
    .C(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__clkbuf_8 _11383_ (.A(net224),
    .X(_06428_));
 sky130_fd_sc_hd__and2_4 _11384_ (.A(_06347_),
    .B(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__a32o_1 _11385_ (.A1(\cur_mb_mem[201][7] ),
    .A2(_06336_),
    .A3(_06093_),
    .B1(_06429_),
    .B2(\cur_mb_mem[67][7] ),
    .X(_06430_));
 sky130_fd_sc_hd__a311o_1 _11386_ (.A1(\cur_mb_mem[249][7] ),
    .A2(_04432_),
    .A3(_05912_),
    .B1(_06427_),
    .C1(_06430_),
    .X(_06431_));
 sky130_fd_sc_hd__and2_4 _11387_ (.A(_05896_),
    .B(_06053_),
    .X(_06432_));
 sky130_fd_sc_hd__and2_4 _11388_ (.A(_05979_),
    .B(_05971_),
    .X(_06433_));
 sky130_fd_sc_hd__clkbuf_8 _11389_ (.A(_05977_),
    .X(_06434_));
 sky130_fd_sc_hd__buf_8 _11390_ (.A(_05953_),
    .X(_06435_));
 sky130_fd_sc_hd__and2_4 _11391_ (.A(_06434_),
    .B(_06435_),
    .X(_06436_));
 sky130_fd_sc_hd__a32o_1 _11392_ (.A1(\cur_mb_mem[173][7] ),
    .A2(_05961_),
    .A3(_06426_),
    .B1(_06436_),
    .B2(\cur_mb_mem[158][7] ),
    .X(_06437_));
 sky130_fd_sc_hd__a221o_1 _11393_ (.A1(\cur_mb_mem[120][7] ),
    .A2(_06432_),
    .B1(_06433_),
    .B2(\cur_mb_mem[144][7] ),
    .C1(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__and2_4 _11394_ (.A(_06051_),
    .B(_06009_),
    .X(_06439_));
 sky130_fd_sc_hd__and2_1 _11395_ (.A(_05904_),
    .B(net225),
    .X(_06440_));
 sky130_fd_sc_hd__clkbuf_16 _11396_ (.A(_06440_),
    .X(_06441_));
 sky130_fd_sc_hd__clkbuf_16 _11397_ (.A(_05903_),
    .X(_06442_));
 sky130_fd_sc_hd__and2_4 _11398_ (.A(_06032_),
    .B(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__a32o_1 _11399_ (.A1(\cur_mb_mem[60][7] ),
    .A2(_05058_),
    .A3(_05989_),
    .B1(_06443_),
    .B2(\cur_mb_mem[250][7] ),
    .X(_06444_));
 sky130_fd_sc_hd__a221o_1 _11400_ (.A1(\cur_mb_mem[112][7] ),
    .A2(_06439_),
    .B1(_06441_),
    .B2(\cur_mb_mem[42][7] ),
    .C1(_06444_),
    .X(_06445_));
 sky130_fd_sc_hd__or4_1 _11401_ (.A(_06425_),
    .B(_06431_),
    .C(_06438_),
    .D(_06445_),
    .X(_06446_));
 sky130_fd_sc_hd__and2_4 _11402_ (.A(_06270_),
    .B(_06179_),
    .X(_06447_));
 sky130_fd_sc_hd__a32o_2 _11403_ (.A1(\cur_mb_mem[222][7] ),
    .A2(_06106_),
    .A3(_06025_),
    .B1(_06447_),
    .B2(\cur_mb_mem[215][7] ),
    .X(_06448_));
 sky130_fd_sc_hd__and2_4 _11404_ (.A(_06442_),
    .B(_06403_),
    .X(_06449_));
 sky130_fd_sc_hd__a32o_1 _11405_ (.A1(\cur_mb_mem[109][7] ),
    .A2(_06298_),
    .A3(_05946_),
    .B1(_06449_),
    .B2(\cur_mb_mem[26][7] ),
    .X(_06450_));
 sky130_fd_sc_hd__and3_1 _11406_ (.A(\cur_mb_mem[192][7] ),
    .B(_06092_),
    .C(_05971_),
    .X(_06451_));
 sky130_fd_sc_hd__a31o_1 _11407_ (.A1(\cur_mb_mem[175][7] ),
    .A2(_04424_),
    .A3(_05923_),
    .B1(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__and2_4 _11408_ (.A(_05909_),
    .B(_06188_),
    .X(_06453_));
 sky130_fd_sc_hd__a32o_1 _11409_ (.A1(\cur_mb_mem[81][7] ),
    .A2(_05925_),
    .A3(_05994_),
    .B1(_06453_),
    .B2(\cur_mb_mem[153][7] ),
    .X(_06454_));
 sky130_fd_sc_hd__buf_12 _11410_ (.A(net255),
    .X(_06455_));
 sky130_fd_sc_hd__clkbuf_8 _11411_ (.A(_06081_),
    .X(_06456_));
 sky130_fd_sc_hd__and2_4 _11412_ (.A(_06455_),
    .B(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__a32o_1 _11413_ (.A1(\cur_mb_mem[168][7] ),
    .A2(_05896_),
    .A3(_06426_),
    .B1(_06457_),
    .B2(\cur_mb_mem[200][7] ),
    .X(_06458_));
 sky130_fd_sc_hd__or4_1 _11414_ (.A(_06450_),
    .B(_06452_),
    .C(_06454_),
    .D(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__and2_4 _11415_ (.A(_06233_),
    .B(_06179_),
    .X(_06460_));
 sky130_fd_sc_hd__buf_12 _11416_ (.A(_06095_),
    .X(_06461_));
 sky130_fd_sc_hd__and2_4 _11417_ (.A(_06461_),
    .B(_05933_),
    .X(_06462_));
 sky130_fd_sc_hd__and2_4 _11418_ (.A(_05896_),
    .B(_06224_),
    .X(_06463_));
 sky130_fd_sc_hd__a32o_1 _11419_ (.A1(\cur_mb_mem[113][7] ),
    .A2(_06119_),
    .A3(_05994_),
    .B1(_06463_),
    .B2(\cur_mb_mem[232][7] ),
    .X(_06464_));
 sky130_fd_sc_hd__a221o_2 _11420_ (.A1(\cur_mb_mem[71][7] ),
    .A2(_06460_),
    .B1(_06462_),
    .B2(\cur_mb_mem[135][7] ),
    .C1(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__buf_8 _11421_ (.A(_06099_),
    .X(_06466_));
 sky130_fd_sc_hd__and2_2 _11422_ (.A(_06466_),
    .B(_06019_),
    .X(_06467_));
 sky130_fd_sc_hd__a32o_2 _11423_ (.A1(\cur_mb_mem[87][7] ),
    .A2(_05916_),
    .A3(_06103_),
    .B1(_06467_),
    .B2(\cur_mb_mem[191][7] ),
    .X(_06468_));
 sky130_fd_sc_hd__or4_1 _11424_ (.A(_06448_),
    .B(_06459_),
    .C(_06465_),
    .D(_06468_),
    .X(_06469_));
 sky130_fd_sc_hd__and3_1 _11425_ (.A(\cur_mb_mem[126][7] ),
    .B(_06118_),
    .C(_05954_),
    .X(_06470_));
 sky130_fd_sc_hd__a31o_1 _11426_ (.A1(\cur_mb_mem[187][7] ),
    .A2(_05919_),
    .A3(_06037_),
    .B1(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__and3_1 _11427_ (.A(\cur_mb_mem[115][7] ),
    .B(_06063_),
    .C(_06118_),
    .X(_06472_));
 sky130_fd_sc_hd__a31o_1 _11428_ (.A1(\cur_mb_mem[169][7] ),
    .A2(_05911_),
    .A3(_06426_),
    .B1(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__buf_12 _11429_ (.A(_05917_),
    .X(_06474_));
 sky130_fd_sc_hd__buf_8 _11430_ (.A(net232),
    .X(_06475_));
 sky130_fd_sc_hd__and2_4 _11431_ (.A(_06474_),
    .B(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__a32o_1 _11432_ (.A1(\cur_mb_mem[195][7] ),
    .A2(_06063_),
    .A3(_06093_),
    .B1(_06476_),
    .B2(\cur_mb_mem[27][7] ),
    .X(_06477_));
 sky130_fd_sc_hd__buf_12 _11433_ (.A(net259),
    .X(_06478_));
 sky130_fd_sc_hd__and2_4 _11434_ (.A(_06478_),
    .B(_06019_),
    .X(_06479_));
 sky130_fd_sc_hd__and2_4 _11435_ (.A(_06039_),
    .B(_06046_),
    .X(_06480_));
 sky130_fd_sc_hd__a22o_1 _11436_ (.A1(\cur_mb_mem[184][7] ),
    .A2(_06479_),
    .B1(_06480_),
    .B2(\cur_mb_mem[190][7] ),
    .X(_06481_));
 sky130_fd_sc_hd__or4_2 _11437_ (.A(_06471_),
    .B(_06473_),
    .C(_06477_),
    .D(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__and2_4 _11438_ (.A(_06428_),
    .B(_06076_),
    .X(_06483_));
 sky130_fd_sc_hd__a32o_1 _11439_ (.A1(\cur_mb_mem[58][7] ),
    .A2(_05059_),
    .A3(_06035_),
    .B1(_06483_),
    .B2(\cur_mb_mem[65][7] ),
    .X(_06484_));
 sky130_fd_sc_hd__nor2_8 _11440_ (.A(_06276_),
    .B(_06258_),
    .Y(_06485_));
 sky130_fd_sc_hd__a32o_1 _11441_ (.A1(\cur_mb_mem[204][7] ),
    .A2(_05989_),
    .A3(_06094_),
    .B1(_06485_),
    .B2(\cur_mb_mem[40][7] ),
    .X(_06486_));
 sky130_fd_sc_hd__and2_4 _11442_ (.A(_06435_),
    .B(_06382_),
    .X(_06487_));
 sky130_fd_sc_hd__buf_4 _11443_ (.A(net232),
    .X(_06488_));
 sky130_fd_sc_hd__and2_4 _11444_ (.A(_06327_),
    .B(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__buf_6 _11445_ (.A(_05944_),
    .X(_06490_));
 sky130_fd_sc_hd__and2_4 _11446_ (.A(_06343_),
    .B(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__a32o_1 _11447_ (.A1(\cur_mb_mem[106][7] ),
    .A2(_06035_),
    .A3(_06299_),
    .B1(_06491_),
    .B2(\cur_mb_mem[45][7] ),
    .X(_06492_));
 sky130_fd_sc_hd__a221o_2 _11448_ (.A1(\cur_mb_mem[142][7] ),
    .A2(_06487_),
    .B1(_06489_),
    .B2(\cur_mb_mem[25][7] ),
    .C1(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__or4_1 _11449_ (.A(_06482_),
    .B(_06484_),
    .C(_06486_),
    .D(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__or4_2 _11450_ (.A(_06420_),
    .B(_06446_),
    .C(_06469_),
    .D(_06494_),
    .X(_06495_));
 sky130_fd_sc_hd__or4_4 _11451_ (.A(_06320_),
    .B(_06332_),
    .C(_06392_),
    .D(_06495_),
    .X(_06496_));
 sky130_fd_sc_hd__o22ai_2 _11452_ (.A1(\cur_mb_mem[0][7] ),
    .A2(_05908_),
    .B1(_06311_),
    .B2(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__nor2_2 _11453_ (.A(net104),
    .B(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__a22o_1 _11454_ (.A1(\cur_mb_mem[162][6] ),
    .A2(_06284_),
    .B1(_06028_),
    .B2(\cur_mb_mem[100][6] ),
    .X(_06499_));
 sky130_fd_sc_hd__a32o_4 _11455_ (.A1(\cur_mb_mem[227][6] ),
    .A2(_06064_),
    .A3(_06067_),
    .B1(_06114_),
    .B2(\cur_mb_mem[7][6] ),
    .X(_06500_));
 sky130_fd_sc_hd__a221o_1 _11456_ (.A1(\cur_mb_mem[74][6] ),
    .A2(_06417_),
    .B1(_06122_),
    .B2(\cur_mb_mem[79][6] ),
    .C1(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__a32o_1 _11457_ (.A1(\cur_mb_mem[198][6] ),
    .A2(_06187_),
    .A3(_06094_),
    .B1(_06148_),
    .B2(\cur_mb_mem[133][6] ),
    .X(_06502_));
 sky130_fd_sc_hd__a32o_1 _11458_ (.A1(\cur_mb_mem[60][6] ),
    .A2(_05059_),
    .A3(_05989_),
    .B1(_06432_),
    .B2(\cur_mb_mem[120][6] ),
    .X(_06503_));
 sky130_fd_sc_hd__a32o_1 _11459_ (.A1(\cur_mb_mem[175][6] ),
    .A2(_04424_),
    .A3(_06426_),
    .B1(_06295_),
    .B2(\cur_mb_mem[15][6] ),
    .X(_06504_));
 sky130_fd_sc_hd__a32o_1 _11460_ (.A1(\cur_mb_mem[109][6] ),
    .A2(_06299_),
    .A3(_05961_),
    .B1(_06305_),
    .B2(\cur_mb_mem[143][6] ),
    .X(_06505_));
 sky130_fd_sc_hd__a22o_1 _11461_ (.A1(\cur_mb_mem[98][6] ),
    .A2(_06330_),
    .B1(_06483_),
    .B2(\cur_mb_mem[65][6] ),
    .X(_06506_));
 sky130_fd_sc_hd__a221o_1 _11462_ (.A1(\cur_mb_mem[101][6] ),
    .A2(_06269_),
    .B1(_06404_),
    .B2(\cur_mb_mem[29][6] ),
    .C1(_06506_),
    .X(_06507_));
 sky130_fd_sc_hd__and3_1 _11463_ (.A(\cur_mb_mem[59][6] ),
    .B(_05057_),
    .C(_05919_),
    .X(_06508_));
 sky130_fd_sc_hd__a32o_1 _11464_ (.A1(\cur_mb_mem[64][6] ),
    .A2(_06024_),
    .A3(_05971_),
    .B1(_06342_),
    .B2(\cur_mb_mem[210][6] ),
    .X(_06509_));
 sky130_fd_sc_hd__a311o_2 _11465_ (.A1(\cur_mb_mem[217][6] ),
    .A2(_06336_),
    .A3(_05942_),
    .B1(_06508_),
    .C1(_06509_),
    .X(_06510_));
 sky130_fd_sc_hd__or4_1 _11466_ (.A(_06504_),
    .B(_06505_),
    .C(_06507_),
    .D(_06510_),
    .X(_06511_));
 sky130_fd_sc_hd__a2111o_1 _11467_ (.A1(\cur_mb_mem[95][6] ),
    .A2(_06297_),
    .B1(_06502_),
    .C1(_06503_),
    .D1(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__a2111o_1 _11468_ (.A1(\cur_mb_mem[31][6] ),
    .A2(_06178_),
    .B1(_06499_),
    .C1(_06501_),
    .D1(_06512_),
    .X(_06513_));
 sky130_fd_sc_hd__a221o_2 _11469_ (.A1(\cur_mb_mem[223][6] ),
    .A2(_06151_),
    .B1(_06174_),
    .B2(\cur_mb_mem[159][6] ),
    .C1(_06513_),
    .X(_06514_));
 sky130_fd_sc_hd__a32o_1 _11470_ (.A1(\cur_mb_mem[48][6] ),
    .A2(_05057_),
    .A3(_05972_),
    .B1(_06075_),
    .B2(\cur_mb_mem[128][6] ),
    .X(_06515_));
 sky130_fd_sc_hd__a221o_1 _11471_ (.A1(\cur_mb_mem[138][6] ),
    .A2(_05934_),
    .B1(_05998_),
    .B2(\cur_mb_mem[225][6] ),
    .C1(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__and3_1 _11472_ (.A(\cur_mb_mem[235][6] ),
    .B(_06261_),
    .C(_06224_),
    .X(_06517_));
 sky130_fd_sc_hd__a31o_1 _11473_ (.A1(\cur_mb_mem[201][6] ),
    .A2(_05911_),
    .A3(_06093_),
    .B1(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__a221o_1 _11474_ (.A1(\cur_mb_mem[135][6] ),
    .A2(_06462_),
    .B1(_06180_),
    .B2(\cur_mb_mem[231][6] ),
    .C1(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__a32o_1 _11475_ (.A1(\cur_mb_mem[228][6] ),
    .A2(_06223_),
    .A3(_06066_),
    .B1(_06318_),
    .B2(\cur_mb_mem[17][6] ),
    .X(_06520_));
 sky130_fd_sc_hd__a221o_1 _11476_ (.A1(\cur_mb_mem[39][6] ),
    .A2(_06373_),
    .B1(_06259_),
    .B2(\cur_mb_mem[47][6] ),
    .C1(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__a32o_1 _11477_ (.A1(\cur_mb_mem[157][6] ),
    .A2(_05946_),
    .A3(_05979_),
    .B1(_06205_),
    .B2(\cur_mb_mem[182][6] ),
    .X(_06522_));
 sky130_fd_sc_hd__a221o_1 _11478_ (.A1(\cur_mb_mem[37][6] ),
    .A2(_06344_),
    .B1(_06189_),
    .B2(\cur_mb_mem[150][6] ),
    .C1(_06522_),
    .X(_06523_));
 sky130_fd_sc_hd__or4_1 _11479_ (.A(_06516_),
    .B(_06519_),
    .C(_06521_),
    .D(_06523_),
    .X(_06524_));
 sky130_fd_sc_hd__a32o_1 _11480_ (.A1(\cur_mb_mem[240][6] ),
    .A2(_04431_),
    .A3(_05973_),
    .B1(_06162_),
    .B2(\cur_mb_mem[4][6] ),
    .X(_06525_));
 sky130_fd_sc_hd__and3_1 _11481_ (.A(\cur_mb_mem[147][6] ),
    .B(_06063_),
    .C(_05979_),
    .X(_06526_));
 sky130_fd_sc_hd__a31o_1 _11482_ (.A1(\cur_mb_mem[252][6] ),
    .A2(_04431_),
    .A3(_05989_),
    .B1(_06526_),
    .X(_06527_));
 sky130_fd_sc_hd__and3_1 _11483_ (.A(\cur_mb_mem[126][6] ),
    .B(_06053_),
    .C(_05955_),
    .X(_06528_));
 sky130_fd_sc_hd__a32o_1 _11484_ (.A1(\cur_mb_mem[32][6] ),
    .A2(_06044_),
    .A3(_05972_),
    .B1(_06393_),
    .B2(\cur_mb_mem[34][6] ),
    .X(_06529_));
 sky130_fd_sc_hd__a311o_1 _11485_ (.A1(\cur_mb_mem[249][6] ),
    .A2(_04431_),
    .A3(_06336_),
    .B1(_06528_),
    .C1(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__a32o_1 _11486_ (.A1(\cur_mb_mem[171][6] ),
    .A2(_05919_),
    .A3(_06137_),
    .B1(_06443_),
    .B2(\cur_mb_mem[250][6] ),
    .X(_06531_));
 sky130_fd_sc_hd__a32o_1 _11487_ (.A1(\cur_mb_mem[90][6] ),
    .A2(_05958_),
    .A3(_05915_),
    .B1(_06034_),
    .B2(\cur_mb_mem[253][6] ),
    .X(_06532_));
 sky130_fd_sc_hd__a32o_2 _11488_ (.A1(\cur_mb_mem[81][6] ),
    .A2(_05915_),
    .A3(_05993_),
    .B1(_06002_),
    .B2(\cur_mb_mem[30][6] ),
    .X(_06533_));
 sky130_fd_sc_hd__a32o_1 _11489_ (.A1(\cur_mb_mem[206][6] ),
    .A2(_05955_),
    .A3(_06093_),
    .B1(_06242_),
    .B2(\cur_mb_mem[22][6] ),
    .X(_06534_));
 sky130_fd_sc_hd__or4_1 _11490_ (.A(_06531_),
    .B(_06532_),
    .C(_06533_),
    .D(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__or4_1 _11491_ (.A(_06525_),
    .B(_06527_),
    .C(_06530_),
    .D(_06535_),
    .X(_06536_));
 sky130_fd_sc_hd__a32o_1 _11492_ (.A1(\cur_mb_mem[113][6] ),
    .A2(_06053_),
    .A3(_05993_),
    .B1(_06335_),
    .B2(\cur_mb_mem[242][6] ),
    .X(_06537_));
 sky130_fd_sc_hd__a221o_1 _11493_ (.A1(\cur_mb_mem[85][6] ),
    .A2(_06231_),
    .B1(_06285_),
    .B2(\cur_mb_mem[24][6] ),
    .C1(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__a32o_1 _11494_ (.A1(\cur_mb_mem[96][6] ),
    .A2(_06298_),
    .A3(_05971_),
    .B1(_06314_),
    .B2(\cur_mb_mem[107][6] ),
    .X(_06539_));
 sky130_fd_sc_hd__a221o_1 _11495_ (.A1(\cur_mb_mem[194][6] ),
    .A2(_06083_),
    .B1(_06088_),
    .B2(\cur_mb_mem[35][6] ),
    .C1(_06539_),
    .X(_06540_));
 sky130_fd_sc_hd__a22o_1 _11496_ (.A1(\cur_mb_mem[132][6] ),
    .A2(net220),
    .B1(_05990_),
    .B2(\cur_mb_mem[1][6] ),
    .X(_06541_));
 sky130_fd_sc_hd__a221o_1 _11497_ (.A1(\cur_mb_mem[52][6] ),
    .A2(_06241_),
    .B1(_06031_),
    .B2(\cur_mb_mem[41][6] ),
    .C1(_06541_),
    .X(_06542_));
 sky130_fd_sc_hd__a32o_1 _11498_ (.A1(\cur_mb_mem[172][6] ),
    .A2(_05937_),
    .A3(_06137_),
    .B1(_06489_),
    .B2(\cur_mb_mem[25][6] ),
    .X(_06543_));
 sky130_fd_sc_hd__a32o_1 _11499_ (.A1(\cur_mb_mem[18][6] ),
    .A2(_06283_),
    .A3(_05976_),
    .B1(\cur_mb_mem[10][6] ),
    .B2(_06408_),
    .X(_06544_));
 sky130_fd_sc_hd__or4_1 _11500_ (.A(_06540_),
    .B(_06542_),
    .C(_06543_),
    .D(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__a32o_1 _11501_ (.A1(\cur_mb_mem[49][6] ),
    .A2(_05057_),
    .A3(_05994_),
    .B1(_06217_),
    .B2(\cur_mb_mem[180][6] ),
    .X(_06546_));
 sky130_fd_sc_hd__a221o_1 _11502_ (.A1(\cur_mb_mem[108][6] ),
    .A2(_06322_),
    .B1(_06291_),
    .B2(\cur_mb_mem[33][6] ),
    .C1(_06546_),
    .X(_06547_));
 sky130_fd_sc_hd__and3_1 _11503_ (.A(\cur_mb_mem[124][6] ),
    .B(_05937_),
    .C(_06052_),
    .X(_06548_));
 sky130_fd_sc_hd__a32o_1 _11504_ (.A1(\cur_mb_mem[154][6] ),
    .A2(_05958_),
    .A3(_05978_),
    .B1(_06441_),
    .B2(\cur_mb_mem[42][6] ),
    .X(_06549_));
 sky130_fd_sc_hd__a311o_4 _11505_ (.A1(\cur_mb_mem[115][6] ),
    .A2(_06063_),
    .A3(_06118_),
    .B1(_06548_),
    .C1(_06549_),
    .X(_06550_));
 sky130_fd_sc_hd__and3_1 _11506_ (.A(\cur_mb_mem[93][6] ),
    .B(_05915_),
    .C(_05945_),
    .X(_06551_));
 sky130_fd_sc_hd__a32o_1 _11507_ (.A1(\cur_mb_mem[51][6] ),
    .A2(_05056_),
    .A3(_06062_),
    .B1(_06356_),
    .B2(\cur_mb_mem[179][6] ),
    .X(_06552_));
 sky130_fd_sc_hd__a311o_1 _11508_ (.A1(\cur_mb_mem[75][6] ),
    .A2(_05919_),
    .A3(_06024_),
    .B1(_06551_),
    .C1(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__a32o_1 _11509_ (.A1(\cur_mb_mem[165][6] ),
    .A2(_05923_),
    .A3(_06133_),
    .B1(\cur_mb_mem[45][6] ),
    .B2(_06491_),
    .X(_06554_));
 sky130_fd_sc_hd__a32o_1 _11510_ (.A1(\cur_mb_mem[160][6] ),
    .A2(_05923_),
    .A3(_05972_),
    .B1(_06351_),
    .B2(\cur_mb_mem[56][6] ),
    .X(_06555_));
 sky130_fd_sc_hd__or4_1 _11511_ (.A(_06550_),
    .B(_06553_),
    .C(_06554_),
    .D(_06555_),
    .X(_06556_));
 sky130_fd_sc_hd__or4_2 _11512_ (.A(_06538_),
    .B(_06545_),
    .C(_06547_),
    .D(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__or3_1 _11513_ (.A(_06524_),
    .B(_06536_),
    .C(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__a32o_1 _11514_ (.A1(\cur_mb_mem[103][6] ),
    .A2(_06299_),
    .A3(_06098_),
    .B1(_06256_),
    .B2(\cur_mb_mem[226][6] ),
    .X(_06559_));
 sky130_fd_sc_hd__a32o_1 _11515_ (.A1(\cur_mb_mem[230][6] ),
    .A2(_06187_),
    .A3(_06067_),
    .B1(_06467_),
    .B2(\cur_mb_mem[191][6] ),
    .X(_06560_));
 sky130_fd_sc_hd__a211o_1 _11516_ (.A1(\cur_mb_mem[127][6] ),
    .A2(_06101_),
    .B1(_06559_),
    .C1(_06560_),
    .X(_06561_));
 sky130_fd_sc_hd__and3_1 _11517_ (.A(\cur_mb_mem[183][6] ),
    .B(_06037_),
    .C(_06097_),
    .X(_06562_));
 sky130_fd_sc_hd__a31o_1 _11518_ (.A1(\cur_mb_mem[87][6] ),
    .A2(_05916_),
    .A3(_06098_),
    .B1(_06562_),
    .X(_06563_));
 sky130_fd_sc_hd__a32o_1 _11519_ (.A1(\cur_mb_mem[238][6] ),
    .A2(_05955_),
    .A3(_06066_),
    .B1(_06069_),
    .B2(\cur_mb_mem[111][6] ),
    .X(_06564_));
 sky130_fd_sc_hd__and3_1 _11520_ (.A(\cur_mb_mem[55][6] ),
    .B(_05056_),
    .C(_06096_),
    .X(_06565_));
 sky130_fd_sc_hd__a31o_1 _11521_ (.A1(\cur_mb_mem[119][6] ),
    .A2(_06118_),
    .A3(_06097_),
    .B1(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__a32o_1 _11522_ (.A1(\cur_mb_mem[63][6] ),
    .A2(_04424_),
    .A3(_05057_),
    .B1(_06304_),
    .B2(\cur_mb_mem[255][6] ),
    .X(_06567_));
 sky130_fd_sc_hd__or2_1 _11523_ (.A(_06566_),
    .B(_06567_),
    .X(_06568_));
 sky130_fd_sc_hd__a32o_1 _11524_ (.A1(\cur_mb_mem[233][6] ),
    .A2(_05910_),
    .A3(_06066_),
    .B1(_06125_),
    .B2(\cur_mb_mem[239][6] ),
    .X(_06569_));
 sky130_fd_sc_hd__a32o_1 _11525_ (.A1(\cur_mb_mem[236][6] ),
    .A2(_05937_),
    .A3(_06066_),
    .B1(_06248_),
    .B2(\cur_mb_mem[237][6] ),
    .X(_06570_));
 sky130_fd_sc_hd__a32o_1 _11526_ (.A1(\cur_mb_mem[199][6] ),
    .A2(_06092_),
    .A3(_06097_),
    .B1(_06117_),
    .B2(\cur_mb_mem[234][6] ),
    .X(_06571_));
 sky130_fd_sc_hd__and3_1 _11527_ (.A(\cur_mb_mem[197][6] ),
    .B(_06091_),
    .C(_06132_),
    .X(_06572_));
 sky130_fd_sc_hd__a31o_1 _11528_ (.A1(\cur_mb_mem[221][6] ),
    .A2(_05946_),
    .A3(_05948_),
    .B1(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__or4_1 _11529_ (.A(_06569_),
    .B(_06570_),
    .C(_06571_),
    .D(_06573_),
    .X(_06574_));
 sky130_fd_sc_hd__or4_1 _11530_ (.A(_06563_),
    .B(_06564_),
    .C(_06568_),
    .D(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__a32o_1 _11531_ (.A1(\cur_mb_mem[208][6] ),
    .A2(_06106_),
    .A3(_05973_),
    .B1(_06325_),
    .B2(\cur_mb_mem[203][6] ),
    .X(_06576_));
 sky130_fd_sc_hd__a32o_4 _11532_ (.A1(\cur_mb_mem[106][6] ),
    .A2(_06035_),
    .A3(_06299_),
    .B1(_06010_),
    .B2(\cur_mb_mem[80][6] ),
    .X(_06577_));
 sky130_fd_sc_hd__and3_1 _11533_ (.A(\cur_mb_mem[170][6] ),
    .B(_05959_),
    .C(_05923_),
    .X(_06578_));
 sky130_fd_sc_hd__a32o_1 _11534_ (.A1(\cur_mb_mem[99][6] ),
    .A2(_06298_),
    .A3(_06063_),
    .B1(_06157_),
    .B2(\cur_mb_mem[5][6] ),
    .X(_06579_));
 sky130_fd_sc_hd__a311o_1 _11535_ (.A1(\cur_mb_mem[213][6] ),
    .A2(_06106_),
    .A3(_06133_),
    .B1(_06578_),
    .C1(_06579_),
    .X(_06580_));
 sky130_fd_sc_hd__a32o_1 _11536_ (.A1(\cur_mb_mem[168][6] ),
    .A2(_05896_),
    .A3(_06137_),
    .B1(_06290_),
    .B2(\cur_mb_mem[3][6] ),
    .X(_06581_));
 sky130_fd_sc_hd__a32o_2 _11537_ (.A1(\cur_mb_mem[23][6] ),
    .A2(_06097_),
    .A3(_05976_),
    .B1(_06014_),
    .B2(\cur_mb_mem[189][6] ),
    .X(_06582_));
 sky130_fd_sc_hd__a22o_1 _11538_ (.A1(\cur_mb_mem[130][6] ),
    .A2(_06266_),
    .B1(_05936_),
    .B2(\cur_mb_mem[137][6] ),
    .X(_06583_));
 sky130_fd_sc_hd__a32o_1 _11539_ (.A1(\cur_mb_mem[54][6] ),
    .A2(_05057_),
    .A3(_06187_),
    .B1(_06288_),
    .B2(\cur_mb_mem[72][6] ),
    .X(_06584_));
 sky130_fd_sc_hd__or4_4 _11540_ (.A(_06581_),
    .B(_06582_),
    .C(_06583_),
    .D(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__or4_1 _11541_ (.A(_06576_),
    .B(_06577_),
    .C(_06580_),
    .D(_06585_),
    .X(_06586_));
 sky130_fd_sc_hd__or4_2 _11542_ (.A(_06185_),
    .B(_06561_),
    .C(_06575_),
    .D(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__and3_1 _11543_ (.A(\cur_mb_mem[9][6] ),
    .B(_06112_),
    .C(_05911_),
    .X(_06588_));
 sky130_fd_sc_hd__and3_1 _11544_ (.A(\cur_mb_mem[187][6] ),
    .B(_06261_),
    .C(_06036_),
    .X(_06589_));
 sky130_fd_sc_hd__a31o_1 _11545_ (.A1(\cur_mb_mem[13][6] ),
    .A2(_06112_),
    .A3(_05961_),
    .B1(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__a311o_1 _11546_ (.A1(\cur_mb_mem[220][6] ),
    .A2(_05989_),
    .A3(_06106_),
    .B1(_06588_),
    .C1(_06590_),
    .X(_06591_));
 sky130_fd_sc_hd__a32o_1 _11547_ (.A1(\cur_mb_mem[163][6] ),
    .A2(_06064_),
    .A3(_05956_),
    .B1(_06020_),
    .B2(\cur_mb_mem[177][6] ),
    .X(_06592_));
 sky130_fd_sc_hd__and3_1 _11548_ (.A(\cur_mb_mem[245][6] ),
    .B(_04431_),
    .C(_06133_),
    .X(_06593_));
 sky130_fd_sc_hd__a31o_1 _11549_ (.A1(\cur_mb_mem[254][6] ),
    .A2(_04432_),
    .A3(_05955_),
    .B1(_06593_),
    .X(_06594_));
 sky130_fd_sc_hd__and3_1 _11550_ (.A(\cur_mb_mem[204][6] ),
    .B(_05937_),
    .C(_06092_),
    .X(_06595_));
 sky130_fd_sc_hd__a31o_1 _11551_ (.A1(\cur_mb_mem[94][6] ),
    .A2(_05915_),
    .A3(_05955_),
    .B1(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__a32o_2 _11552_ (.A1(\cur_mb_mem[148][6] ),
    .A2(_06223_),
    .A3(_05979_),
    .B1(_06234_),
    .B2(\cur_mb_mem[68][6] ),
    .X(_06597_));
 sky130_fd_sc_hd__a32o_1 _11553_ (.A1(\cur_mb_mem[243][6] ),
    .A2(_04430_),
    .A3(_06063_),
    .B1(_06399_),
    .B2(\cur_mb_mem[44][6] ),
    .X(_06598_));
 sky130_fd_sc_hd__a22o_1 _11554_ (.A1(\cur_mb_mem[102][6] ),
    .A2(_06414_),
    .B1(_06277_),
    .B2(\cur_mb_mem[8][6] ),
    .X(_06599_));
 sky130_fd_sc_hd__or4_1 _11555_ (.A(_06596_),
    .B(_06597_),
    .C(_06598_),
    .D(_06599_),
    .X(_06600_));
 sky130_fd_sc_hd__or4_1 _11556_ (.A(_06591_),
    .B(_06592_),
    .C(_06594_),
    .D(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__and3_1 _11557_ (.A(\cur_mb_mem[149][6] ),
    .B(_05978_),
    .C(_06132_),
    .X(_06602_));
 sky130_fd_sc_hd__a32o_2 _11558_ (.A1(\cur_mb_mem[169][6] ),
    .A2(_05910_),
    .A3(_05922_),
    .B1(_06328_),
    .B2(\cur_mb_mem[73][6] ),
    .X(_06603_));
 sky130_fd_sc_hd__a311o_1 _11559_ (.A1(\cur_mb_mem[251][6] ),
    .A2(_04430_),
    .A3(_05919_),
    .B1(_06602_),
    .C1(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__a32o_2 _11560_ (.A1(\cur_mb_mem[125][6] ),
    .A2(_05945_),
    .A3(_06052_),
    .B1(_06141_),
    .B2(\cur_mb_mem[118][6] ),
    .X(_06605_));
 sky130_fd_sc_hd__a221o_1 _11561_ (.A1(\cur_mb_mem[166][6] ),
    .A2(_06193_),
    .B1(_06480_),
    .B2(\cur_mb_mem[190][6] ),
    .C1(_06605_),
    .X(_06606_));
 sky130_fd_sc_hd__a32o_2 _11562_ (.A1(\cur_mb_mem[123][6] ),
    .A2(_06261_),
    .A3(_06052_),
    .B1(_06077_),
    .B2(\cur_mb_mem[97][6] ),
    .X(_06607_));
 sky130_fd_sc_hd__a221o_1 _11563_ (.A1(\cur_mb_mem[139][6] ),
    .A2(_06388_),
    .B1(_06301_),
    .B2(\cur_mb_mem[11][6] ),
    .C1(_06607_),
    .X(_06608_));
 sky130_fd_sc_hd__a32o_1 _11564_ (.A1(\cur_mb_mem[222][6] ),
    .A2(_05941_),
    .A3(_05954_),
    .B1(_06354_),
    .B2(\cur_mb_mem[193][6] ),
    .X(_06609_));
 sky130_fd_sc_hd__a221o_1 _11565_ (.A1(\cur_mb_mem[141][6] ),
    .A2(_06250_),
    .B1(_06349_),
    .B2(\cur_mb_mem[211][6] ),
    .C1(_06609_),
    .X(_06610_));
 sky130_fd_sc_hd__or4_2 _11566_ (.A(_06604_),
    .B(_06606_),
    .C(_06608_),
    .D(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__a32o_1 _11567_ (.A1(\cur_mb_mem[88][6] ),
    .A2(_05896_),
    .A3(_05925_),
    .B1(_06292_),
    .B2(\cur_mb_mem[136][6] ),
    .X(_06612_));
 sky130_fd_sc_hd__a221o_1 _11568_ (.A1(\cur_mb_mem[91][6] ),
    .A2(_06361_),
    .B1(_06476_),
    .B2(\cur_mb_mem[27][6] ),
    .C1(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__a32o_1 _11569_ (.A1(\cur_mb_mem[174][6] ),
    .A2(_05955_),
    .A3(_05923_),
    .B1(_06439_),
    .B2(\cur_mb_mem[112][6] ),
    .X(_06614_));
 sky130_fd_sc_hd__a32o_1 _11570_ (.A1(\cur_mb_mem[89][6] ),
    .A2(_05911_),
    .A3(_05915_),
    .B1(_06203_),
    .B2(\cur_mb_mem[6][6] ),
    .X(_06615_));
 sky130_fd_sc_hd__a22o_1 _11571_ (.A1(\cur_mb_mem[200][6] ),
    .A2(_06457_),
    .B1(_06423_),
    .B2(\cur_mb_mem[140][6] ),
    .X(_06616_));
 sky130_fd_sc_hd__a221o_1 _11572_ (.A1(\cur_mb_mem[83][6] ),
    .A2(_06379_),
    .B1(_06236_),
    .B2(\cur_mb_mem[21][6] ),
    .C1(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__a32o_1 _11573_ (.A1(\cur_mb_mem[2][6] ),
    .A2(_06112_),
    .A3(_06283_),
    .B1(_06368_),
    .B2(\cur_mb_mem[66][6] ),
    .X(_06618_));
 sky130_fd_sc_hd__a221o_4 _11574_ (.A1(\cur_mb_mem[129][6] ),
    .A2(_05966_),
    .B1(_06172_),
    .B2(\cur_mb_mem[50][6] ),
    .C1(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__or4_1 _11575_ (.A(_06614_),
    .B(_06615_),
    .C(_06617_),
    .D(_06619_),
    .X(_06620_));
 sky130_fd_sc_hd__a32o_1 _11576_ (.A1(\cur_mb_mem[105][6] ),
    .A2(_05910_),
    .A3(_06298_),
    .B1(_06340_),
    .B2(\cur_mb_mem[76][6] ),
    .X(_06621_));
 sky130_fd_sc_hd__a221o_1 _11577_ (.A1(\cur_mb_mem[216][6] ),
    .A2(_06317_),
    .B1(_06411_),
    .B2(\cur_mb_mem[248][6] ),
    .C1(_06621_),
    .X(_06622_));
 sky130_fd_sc_hd__a22o_1 _11578_ (.A1(\cur_mb_mem[146][6] ),
    .A2(_06381_),
    .B1(_06047_),
    .B2(\cur_mb_mem[110][6] ),
    .X(_06623_));
 sky130_fd_sc_hd__a221o_2 _11579_ (.A1(\cur_mb_mem[61][6] ),
    .A2(_06359_),
    .B1(_06239_),
    .B2(\cur_mb_mem[116][6] ),
    .C1(_06623_),
    .X(_06624_));
 sky130_fd_sc_hd__a32o_4 _11580_ (.A1(\cur_mb_mem[122][6] ),
    .A2(_05958_),
    .A3(_06052_),
    .B1(_06370_),
    .B2(\cur_mb_mem[205][6] ),
    .X(_06625_));
 sky130_fd_sc_hd__a221o_1 _11581_ (.A1(\cur_mb_mem[134][6] ),
    .A2(_06211_),
    .B1(_06383_),
    .B2(\cur_mb_mem[131][6] ),
    .C1(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__a32o_4 _11582_ (.A1(\cur_mb_mem[173][6] ),
    .A2(_05945_),
    .A3(_06137_),
    .B1(_06487_),
    .B2(\cur_mb_mem[142][6] ),
    .X(_06627_));
 sky130_fd_sc_hd__a221o_2 _11583_ (.A1(\cur_mb_mem[26][6] ),
    .A2(_06449_),
    .B1(_06017_),
    .B2(\cur_mb_mem[28][6] ),
    .C1(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__or4_1 _11584_ (.A(_06622_),
    .B(_06624_),
    .C(_06626_),
    .D(_06628_),
    .X(_06629_));
 sky130_fd_sc_hd__or4_1 _11585_ (.A(_06611_),
    .B(_06613_),
    .C(_06620_),
    .D(_06629_),
    .X(_06630_));
 sky130_fd_sc_hd__or2_1 _11586_ (.A(_06601_),
    .B(_06630_),
    .X(_06631_));
 sky130_fd_sc_hd__a32o_1 _11587_ (.A1(\cur_mb_mem[229][6] ),
    .A2(_06133_),
    .A3(_06067_),
    .B1(_06460_),
    .B2(\cur_mb_mem[71][6] ),
    .X(_06632_));
 sky130_fd_sc_hd__a221o_1 _11588_ (.A1(\cur_mb_mem[178][6] ),
    .A2(_06386_),
    .B1(_06144_),
    .B2(\cur_mb_mem[70][6] ),
    .C1(_06632_),
    .X(_06633_));
 sky130_fd_sc_hd__and3_1 _11589_ (.A(\cur_mb_mem[224][6] ),
    .B(_05972_),
    .C(_06066_),
    .X(_06634_));
 sky130_fd_sc_hd__a31o_1 _11590_ (.A1(\cur_mb_mem[167][6] ),
    .A2(_05956_),
    .A3(_06098_),
    .B1(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__and3_1 _11591_ (.A(\cur_mb_mem[92][6] ),
    .B(_05938_),
    .C(_05925_),
    .X(_06636_));
 sky130_fd_sc_hd__a31o_1 _11592_ (.A1(\cur_mb_mem[151][6] ),
    .A2(_05980_),
    .A3(_06098_),
    .B1(_06636_),
    .X(_06637_));
 sky130_fd_sc_hd__a32o_1 _11593_ (.A1(\cur_mb_mem[207][6] ),
    .A2(_04424_),
    .A3(_06093_),
    .B1(_06485_),
    .B2(\cur_mb_mem[40][6] ),
    .X(_06638_));
 sky130_fd_sc_hd__a221o_1 _11594_ (.A1(\cur_mb_mem[46][6] ),
    .A2(_06107_),
    .B1(_06433_),
    .B2(\cur_mb_mem[144][6] ),
    .C1(_06638_),
    .X(_06639_));
 sky130_fd_sc_hd__a32o_2 _11595_ (.A1(\cur_mb_mem[247][6] ),
    .A2(_04430_),
    .A3(_06097_),
    .B1(_06463_),
    .B2(\cur_mb_mem[232][6] ),
    .X(_06640_));
 sky130_fd_sc_hd__a221o_2 _11596_ (.A1(\cur_mb_mem[215][6] ),
    .A2(_06447_),
    .B1(_06453_),
    .B2(\cur_mb_mem[153][6] ),
    .C1(_06640_),
    .X(_06641_));
 sky130_fd_sc_hd__or4_1 _11597_ (.A(_06635_),
    .B(_06637_),
    .C(_06639_),
    .D(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__and3_1 _11598_ (.A(\cur_mb_mem[188][6] ),
    .B(_05938_),
    .C(_06037_),
    .X(_06643_));
 sky130_fd_sc_hd__a31o_1 _11599_ (.A1(\cur_mb_mem[121][6] ),
    .A2(_05912_),
    .A3(_06119_),
    .B1(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__a32o_1 _11600_ (.A1(\cur_mb_mem[241][6] ),
    .A2(_04432_),
    .A3(_05994_),
    .B1(_06167_),
    .B2(\cur_mb_mem[244][6] ),
    .X(_06645_));
 sky130_fd_sc_hd__a32o_1 _11601_ (.A1(\cur_mb_mem[86][6] ),
    .A2(_05915_),
    .A3(_06186_),
    .B1(_06280_),
    .B2(\cur_mb_mem[114][6] ),
    .X(_06646_));
 sky130_fd_sc_hd__a221o_1 _11602_ (.A1(\cur_mb_mem[38][6] ),
    .A2(_06396_),
    .B1(_06271_),
    .B2(\cur_mb_mem[209][6] ),
    .C1(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__and3_1 _11603_ (.A(\cur_mb_mem[78][6] ),
    .B(_06023_),
    .C(_05954_),
    .X(_06648_));
 sky130_fd_sc_hd__a31o_1 _11604_ (.A1(\cur_mb_mem[192][6] ),
    .A2(_06093_),
    .A3(_05972_),
    .B1(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__a32o_1 _11605_ (.A1(\cur_mb_mem[202][6] ),
    .A2(_05959_),
    .A3(_06092_),
    .B1(_06334_),
    .B2(\cur_mb_mem[161][6] ),
    .X(_06650_));
 sky130_fd_sc_hd__a32o_1 _11606_ (.A1(\cur_mb_mem[218][6] ),
    .A2(_05958_),
    .A3(_05941_),
    .B1(_06058_),
    .B2(\cur_mb_mem[77][6] ),
    .X(_06651_));
 sky130_fd_sc_hd__a221o_1 _11607_ (.A1(\cur_mb_mem[184][6] ),
    .A2(_06479_),
    .B1(_06218_),
    .B2(\cur_mb_mem[69][6] ),
    .C1(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__or4_1 _11608_ (.A(_06647_),
    .B(_06649_),
    .C(_06650_),
    .D(_06652_),
    .X(_06653_));
 sky130_fd_sc_hd__or3_1 _11609_ (.A(_06644_),
    .B(_06645_),
    .C(_06653_),
    .X(_06654_));
 sky130_fd_sc_hd__and3_1 _11610_ (.A(\cur_mb_mem[20][6] ),
    .B(_06134_),
    .C(_05975_),
    .X(_06655_));
 sky130_fd_sc_hd__a31o_1 _11611_ (.A1(\cur_mb_mem[57][6] ),
    .A2(_05058_),
    .A3(_05911_),
    .B1(_06655_),
    .X(_06656_));
 sky130_fd_sc_hd__a221o_1 _11612_ (.A1(\cur_mb_mem[164][6] ),
    .A2(_06195_),
    .B1(_06402_),
    .B2(\cur_mb_mem[155][6] ),
    .C1(_06656_),
    .X(_06657_));
 sky130_fd_sc_hd__a32o_1 _11613_ (.A1(\cur_mb_mem[62][6] ),
    .A2(_05057_),
    .A3(_05955_),
    .B1(_06135_),
    .B2(\cur_mb_mem[212][6] ),
    .X(_06658_));
 sky130_fd_sc_hd__a32o_1 _11614_ (.A1(\cur_mb_mem[219][6] ),
    .A2(_05919_),
    .A3(_05942_),
    .B1(_06282_),
    .B2(\cur_mb_mem[19][6] ),
    .X(_06659_));
 sky130_fd_sc_hd__a32o_1 _11615_ (.A1(\cur_mb_mem[196][6] ),
    .A2(_05890_),
    .A3(_06091_),
    .B1(_06006_),
    .B2(\cur_mb_mem[43][6] ),
    .X(_06660_));
 sky130_fd_sc_hd__a221o_1 _11616_ (.A1(\cur_mb_mem[36][6] ),
    .A2(_06360_),
    .B1(_06252_),
    .B2(\cur_mb_mem[145][6] ),
    .C1(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__and3_1 _11617_ (.A(\cur_mb_mem[214][6] ),
    .B(_06191_),
    .C(_05947_),
    .X(_06662_));
 sky130_fd_sc_hd__a31o_1 _11618_ (.A1(\cur_mb_mem[84][6] ),
    .A2(_06134_),
    .A3(_05915_),
    .B1(_06662_),
    .X(_06663_));
 sky130_fd_sc_hd__a221o_1 _11619_ (.A1(\cur_mb_mem[117][6] ),
    .A2(_06209_),
    .B1(_06367_),
    .B2(\cur_mb_mem[14][6] ),
    .C1(_06663_),
    .X(_06664_));
 sky130_fd_sc_hd__or4_1 _11620_ (.A(_06658_),
    .B(_06659_),
    .C(_06661_),
    .D(_06664_),
    .X(_06665_));
 sky130_fd_sc_hd__a32o_2 _11621_ (.A1(\cur_mb_mem[156][6] ),
    .A2(_05938_),
    .A3(_05979_),
    .B1(_05985_),
    .B2(\cur_mb_mem[104][6] ),
    .X(_06666_));
 sky130_fd_sc_hd__and3_1 _11622_ (.A(\cur_mb_mem[195][6] ),
    .B(_06062_),
    .C(_06092_),
    .X(_06667_));
 sky130_fd_sc_hd__a31o_1 _11623_ (.A1(\cur_mb_mem[58][6] ),
    .A2(_05057_),
    .A3(_05959_),
    .B1(_06667_),
    .X(_06668_));
 sky130_fd_sc_hd__a32o_1 _11624_ (.A1(\cur_mb_mem[82][6] ),
    .A2(_06283_),
    .A3(_05915_),
    .B1(_06429_),
    .B2(\cur_mb_mem[67][6] ),
    .X(_06669_));
 sky130_fd_sc_hd__a221o_4 _11625_ (.A1(\cur_mb_mem[53][6] ),
    .A2(_06221_),
    .B1(_06316_),
    .B2(\cur_mb_mem[176][6] ),
    .C1(_06669_),
    .X(_06670_));
 sky130_fd_sc_hd__a32o_1 _11626_ (.A1(\cur_mb_mem[181][6] ),
    .A2(_06036_),
    .A3(_06132_),
    .B1(_06160_),
    .B2(\cur_mb_mem[246][6] ),
    .X(_06671_));
 sky130_fd_sc_hd__a32o_1 _11627_ (.A1(\cur_mb_mem[16][6] ),
    .A2(_06315_),
    .A3(_05975_),
    .B1(_06394_),
    .B2(\cur_mb_mem[152][6] ),
    .X(_06672_));
 sky130_fd_sc_hd__a32o_1 _11628_ (.A1(\cur_mb_mem[186][6] ),
    .A2(_05905_),
    .A3(_06036_),
    .B1(_06040_),
    .B2(\cur_mb_mem[185][6] ),
    .X(_06673_));
 sky130_fd_sc_hd__a22o_1 _11629_ (.A1(\cur_mb_mem[12][6] ),
    .A2(_05928_),
    .B1(_06436_),
    .B2(\cur_mb_mem[158][6] ),
    .X(_06674_));
 sky130_fd_sc_hd__or4_1 _11630_ (.A(_06671_),
    .B(_06672_),
    .C(_06673_),
    .D(_06674_),
    .X(_06675_));
 sky130_fd_sc_hd__or4_1 _11631_ (.A(_06666_),
    .B(_06668_),
    .C(_06670_),
    .D(_06675_),
    .X(_06676_));
 sky130_fd_sc_hd__or3_1 _11632_ (.A(_06657_),
    .B(_06665_),
    .C(_06676_),
    .X(_06677_));
 sky130_fd_sc_hd__or4_1 _11633_ (.A(_06633_),
    .B(_06642_),
    .C(_06654_),
    .D(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__or4_4 _11634_ (.A(_06558_),
    .B(_06587_),
    .C(_06631_),
    .D(_06678_),
    .X(_06679_));
 sky130_fd_sc_hd__inv_2 _11635_ (.A(net103),
    .Y(_06680_));
 sky130_fd_sc_hd__o221a_1 _11636_ (.A1(\cur_mb_mem[0][6] ),
    .A2(_05908_),
    .B1(_06514_),
    .B2(_06679_),
    .C1(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__a32o_1 _11637_ (.A1(\cur_mb_mem[123][5] ),
    .A2(_06049_),
    .A3(_06053_),
    .B1(_06394_),
    .B2(\cur_mb_mem[152][5] ),
    .X(_06682_));
 sky130_fd_sc_hd__and3_1 _11638_ (.A(\cur_mb_mem[125][5] ),
    .B(_05945_),
    .C(_06052_),
    .X(_06683_));
 sky130_fd_sc_hd__a31o_1 _11639_ (.A1(\cur_mb_mem[124][5] ),
    .A2(_05938_),
    .A3(_06118_),
    .B1(_06683_),
    .X(_06684_));
 sky130_fd_sc_hd__a32o_1 _11640_ (.A1(\cur_mb_mem[122][5] ),
    .A2(_05959_),
    .A3(_06118_),
    .B1(_06196_),
    .B2(\cur_mb_mem[132][5] ),
    .X(_06685_));
 sky130_fd_sc_hd__a211o_1 _11641_ (.A1(\cur_mb_mem[158][5] ),
    .A2(_06436_),
    .B1(_06684_),
    .C1(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__a211o_1 _11642_ (.A1(\cur_mb_mem[133][5] ),
    .A2(_06148_),
    .B1(_06682_),
    .C1(_06686_),
    .X(_06687_));
 sky130_fd_sc_hd__a32o_1 _11643_ (.A1(\cur_mb_mem[121][5] ),
    .A2(_06336_),
    .A3(_06119_),
    .B1(_06439_),
    .B2(\cur_mb_mem[112][5] ),
    .X(_06688_));
 sky130_fd_sc_hd__a221o_1 _11644_ (.A1(\cur_mb_mem[146][5] ),
    .A2(_06381_),
    .B1(_06231_),
    .B2(\cur_mb_mem[85][5] ),
    .C1(_06688_),
    .X(_06689_));
 sky130_fd_sc_hd__a22o_1 _11645_ (.A1(\cur_mb_mem[118][5] ),
    .A2(_06141_),
    .B1(_06209_),
    .B2(\cur_mb_mem[117][5] ),
    .X(_06690_));
 sky130_fd_sc_hd__a221o_1 _11646_ (.A1(\cur_mb_mem[116][5] ),
    .A2(_06239_),
    .B1(_06402_),
    .B2(\cur_mb_mem[155][5] ),
    .C1(_06690_),
    .X(_06691_));
 sky130_fd_sc_hd__or4_4 _11647_ (.A(_06185_),
    .B(_06687_),
    .C(_06689_),
    .D(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__and3_1 _11648_ (.A(\cur_mb_mem[16][5] ),
    .B(_06074_),
    .C(_06403_),
    .X(_06693_));
 sky130_fd_sc_hd__and3_1 _11649_ (.A(\cur_mb_mem[78][5] ),
    .B(_06143_),
    .C(_06366_),
    .X(_06694_));
 sky130_fd_sc_hd__and3_1 _11650_ (.A(\cur_mb_mem[18][5] ),
    .B(_06341_),
    .C(_06475_),
    .X(_06695_));
 sky130_fd_sc_hd__a2111o_1 _11651_ (.A1(\cur_mb_mem[17][5] ),
    .A2(_06318_),
    .B1(_06693_),
    .C1(_06694_),
    .D1(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__and3_1 _11652_ (.A(\cur_mb_mem[5][5] ),
    .B(_06365_),
    .C(_06131_),
    .X(_06697_));
 sky130_fd_sc_hd__and3_4 _11653_ (.A(\cur_mb_mem[190][5] ),
    .B(_06039_),
    .C(_06366_),
    .X(_06698_));
 sky130_fd_sc_hd__and3_1 _11654_ (.A(\cur_mb_mem[23][5] ),
    .B(_06179_),
    .C(_06475_),
    .X(_06699_));
 sky130_fd_sc_hd__a2111o_1 _11655_ (.A1(\cur_mb_mem[164][5] ),
    .A2(_06195_),
    .B1(_06697_),
    .C1(_06698_),
    .D1(_06699_),
    .X(_06700_));
 sky130_fd_sc_hd__and3_1 _11656_ (.A(\cur_mb_mem[29][5] ),
    .B(_06011_),
    .C(_06403_),
    .X(_06701_));
 sky130_fd_sc_hd__and3_1 _11657_ (.A(\cur_mb_mem[27][5] ),
    .B(_06003_),
    .C(_06488_),
    .X(_06702_));
 sky130_fd_sc_hd__and3_1 _11658_ (.A(\cur_mb_mem[1][5] ),
    .B(_06202_),
    .C(_06353_),
    .X(_06703_));
 sky130_fd_sc_hd__a2111o_1 _11659_ (.A1(\cur_mb_mem[19][5] ),
    .A2(_06282_),
    .B1(_06701_),
    .C1(_06702_),
    .D1(_06703_),
    .X(_06704_));
 sky130_fd_sc_hd__and3_1 _11660_ (.A(\cur_mb_mem[28][5] ),
    .B(_06422_),
    .C(_06475_),
    .X(_06705_));
 sky130_fd_sc_hd__and3_1 _11661_ (.A(\cur_mb_mem[4][5] ),
    .B(_06166_),
    .C(_06300_),
    .X(_06706_));
 sky130_fd_sc_hd__buf_12 _11662_ (.A(net251),
    .X(_06707_));
 sky130_fd_sc_hd__buf_8 _11663_ (.A(_06095_),
    .X(_06708_));
 sky130_fd_sc_hd__and3_1 _11664_ (.A(\cur_mb_mem[7][5] ),
    .B(_06707_),
    .C(_06708_),
    .X(_06709_));
 sky130_fd_sc_hd__a2111o_1 _11665_ (.A1(\cur_mb_mem[12][5] ),
    .A2(_05928_),
    .B1(_06705_),
    .C1(_06706_),
    .D1(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__or4_4 _11666_ (.A(_06696_),
    .B(_06700_),
    .C(_06704_),
    .D(_06710_),
    .X(_06711_));
 sky130_fd_sc_hd__and3_1 _11667_ (.A(\cur_mb_mem[3][5] ),
    .B(_06365_),
    .C(_06061_),
    .X(_06712_));
 sky130_fd_sc_hd__and3_1 _11668_ (.A(\cur_mb_mem[30][5] ),
    .B(_06046_),
    .C(_06488_),
    .X(_06713_));
 sky130_fd_sc_hd__and3_1 _11669_ (.A(\cur_mb_mem[24][5] ),
    .B(_06455_),
    .C(_06475_),
    .X(_06714_));
 sky130_fd_sc_hd__a2111o_1 _11670_ (.A1(\cur_mb_mem[26][5] ),
    .A2(_06449_),
    .B1(_06712_),
    .C1(_06713_),
    .D1(_06714_),
    .X(_06715_));
 sky130_fd_sc_hd__and3_1 _11671_ (.A(\cur_mb_mem[77][5] ),
    .B(_06033_),
    .C(_06428_),
    .X(_06716_));
 sky130_fd_sc_hd__and3_1 _11672_ (.A(\cur_mb_mem[66][5] ),
    .B(_06171_),
    .C(_06143_),
    .X(_06717_));
 sky130_fd_sc_hd__clkbuf_16 _11673_ (.A(_05900_),
    .X(_06718_));
 sky130_fd_sc_hd__and3_1 _11674_ (.A(\cur_mb_mem[76][5] ),
    .B(_06718_),
    .C(_06233_),
    .X(_06719_));
 sky130_fd_sc_hd__a2111o_1 _11675_ (.A1(\cur_mb_mem[72][5] ),
    .A2(_06288_),
    .B1(_06716_),
    .C1(_06717_),
    .D1(_06719_),
    .X(_06720_));
 sky130_fd_sc_hd__and3_1 _11676_ (.A(\cur_mb_mem[22][5] ),
    .B(_06210_),
    .C(_06488_),
    .X(_06721_));
 sky130_fd_sc_hd__and3_1 _11677_ (.A(\cur_mb_mem[75][5] ),
    .B(_06003_),
    .C(_06143_),
    .X(_06722_));
 sky130_fd_sc_hd__buf_8 _11678_ (.A(_05892_),
    .X(_06723_));
 sky130_fd_sc_hd__and3_1 _11679_ (.A(\cur_mb_mem[9][5] ),
    .B(_06202_),
    .C(_06723_),
    .X(_06724_));
 sky130_fd_sc_hd__a2111o_1 _11680_ (.A1(\cur_mb_mem[14][5] ),
    .A2(_06367_),
    .B1(_06721_),
    .C1(_06722_),
    .D1(_06724_),
    .X(_06725_));
 sky130_fd_sc_hd__and3_1 _11681_ (.A(\cur_mb_mem[25][5] ),
    .B(_06327_),
    .C(_06475_),
    .X(_06726_));
 sky130_fd_sc_hd__and3_1 _11682_ (.A(\cur_mb_mem[2][5] ),
    .B(_06202_),
    .C(_06254_),
    .X(_06727_));
 sky130_fd_sc_hd__and3_1 _11683_ (.A(\cur_mb_mem[8][5] ),
    .B(_06707_),
    .C(_05982_),
    .X(_06728_));
 sky130_fd_sc_hd__a2111o_1 _11684_ (.A1(\cur_mb_mem[67][5] ),
    .A2(_06429_),
    .B1(_06726_),
    .C1(_06727_),
    .D1(_06728_),
    .X(_06729_));
 sky130_fd_sc_hd__or4_4 _11685_ (.A(_06715_),
    .B(_06720_),
    .C(_06725_),
    .D(_06729_),
    .X(_06730_));
 sky130_fd_sc_hd__buf_4 _11686_ (.A(_06050_),
    .X(_06731_));
 sky130_fd_sc_hd__and3_1 _11687_ (.A(\cur_mb_mem[113][5] ),
    .B(_06731_),
    .C(_06076_),
    .X(_06732_));
 sky130_fd_sc_hd__and3_1 _11688_ (.A(\cur_mb_mem[114][5] ),
    .B(_06171_),
    .C(_06051_),
    .X(_06733_));
 sky130_fd_sc_hd__and3_1 _11689_ (.A(\cur_mb_mem[119][5] ),
    .B(_06138_),
    .C(_06372_),
    .X(_06734_));
 sky130_fd_sc_hd__a2111o_1 _11690_ (.A1(\cur_mb_mem[43][5] ),
    .A2(_06006_),
    .B1(_06732_),
    .C1(_06733_),
    .D1(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__and3_1 _11691_ (.A(\cur_mb_mem[147][5] ),
    .B(_06347_),
    .C(_06188_),
    .X(_06736_));
 sky130_fd_sc_hd__and3_1 _11692_ (.A(\cur_mb_mem[126][5] ),
    .B(_06051_),
    .C(_06046_),
    .X(_06737_));
 sky130_fd_sc_hd__and3_1 _11693_ (.A(\cur_mb_mem[151][5] ),
    .B(_06401_),
    .C(_06372_),
    .X(_06738_));
 sky130_fd_sc_hd__a2111o_1 _11694_ (.A1(\cur_mb_mem[41][5] ),
    .A2(_06031_),
    .B1(_06736_),
    .C1(_06737_),
    .D1(_06738_),
    .X(_06739_));
 sky130_fd_sc_hd__and3_1 _11695_ (.A(\cur_mb_mem[156][5] ),
    .B(_06422_),
    .C(_06434_),
    .X(_06740_));
 sky130_fd_sc_hd__and3_1 _11696_ (.A(\cur_mb_mem[115][5] ),
    .B(_06355_),
    .C(_06051_),
    .X(_06741_));
 sky130_fd_sc_hd__and3_1 _11697_ (.A(\cur_mb_mem[120][5] ),
    .B(_06478_),
    .C(_06207_),
    .X(_06742_));
 sky130_fd_sc_hd__a2111o_1 _11698_ (.A1(\cur_mb_mem[150][5] ),
    .A2(_06189_),
    .B1(_06740_),
    .C1(_06741_),
    .D1(_06742_),
    .X(_06743_));
 sky130_fd_sc_hd__buf_12 _11699_ (.A(net264),
    .X(_06744_));
 sky130_fd_sc_hd__and3_2 _11700_ (.A(\cur_mb_mem[84][5] ),
    .B(_06744_),
    .C(_06378_),
    .X(_06745_));
 sky130_fd_sc_hd__and3_1 _11701_ (.A(\cur_mb_mem[149][5] ),
    .B(_06401_),
    .C(_06147_),
    .X(_06746_));
 sky130_fd_sc_hd__buf_4 _11702_ (.A(_05977_),
    .X(_06747_));
 sky130_fd_sc_hd__buf_12 _11703_ (.A(net238),
    .X(_06748_));
 sky130_fd_sc_hd__and3_1 _11704_ (.A(\cur_mb_mem[144][5] ),
    .B(_06747_),
    .C(_06748_),
    .X(_06749_));
 sky130_fd_sc_hd__a2111o_1 _11705_ (.A1(\cur_mb_mem[42][5] ),
    .A2(_06441_),
    .B1(_06745_),
    .C1(_06746_),
    .D1(_06749_),
    .X(_06750_));
 sky130_fd_sc_hd__or4_4 _11706_ (.A(_06735_),
    .B(_06739_),
    .C(_06743_),
    .D(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__and3_1 _11707_ (.A(\cur_mb_mem[179][5] ),
    .B(_06355_),
    .C(_06039_),
    .X(_06752_));
 sky130_fd_sc_hd__and3_1 _11708_ (.A(\cur_mb_mem[188][5] ),
    .B(_06718_),
    .C(_06019_),
    .X(_06753_));
 sky130_fd_sc_hd__buf_12 _11709_ (.A(_05900_),
    .X(_06754_));
 sky130_fd_sc_hd__buf_8 _11710_ (.A(_05921_),
    .X(_06755_));
 sky130_fd_sc_hd__and3_1 _11711_ (.A(\cur_mb_mem[172][5] ),
    .B(_06754_),
    .C(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__a2111o_1 _11712_ (.A1(\cur_mb_mem[189][5] ),
    .A2(_06014_),
    .B1(_06752_),
    .C1(_06753_),
    .D1(_06756_),
    .X(_06757_));
 sky130_fd_sc_hd__clkbuf_16 _11713_ (.A(_05920_),
    .X(_06758_));
 sky130_fd_sc_hd__and3_1 _11714_ (.A(\cur_mb_mem[174][5] ),
    .B(_06435_),
    .C(_06758_),
    .X(_06759_));
 sky130_fd_sc_hd__clkbuf_16 _11715_ (.A(_06018_),
    .X(_06760_));
 sky130_fd_sc_hd__and3_1 _11716_ (.A(\cur_mb_mem[187][5] ),
    .B(_06474_),
    .C(_06760_),
    .X(_06761_));
 sky130_fd_sc_hd__buf_8 _11717_ (.A(_05944_),
    .X(_06762_));
 sky130_fd_sc_hd__and3_1 _11718_ (.A(\cur_mb_mem[173][5] ),
    .B(_06762_),
    .C(_06755_),
    .X(_06763_));
 sky130_fd_sc_hd__a2111o_2 _11719_ (.A1(\cur_mb_mem[10][5] ),
    .A2(_06408_),
    .B1(_06759_),
    .C1(_06761_),
    .D1(_06763_),
    .X(_06764_));
 sky130_fd_sc_hd__and3_1 _11720_ (.A(\cur_mb_mem[233][5] ),
    .B(_06327_),
    .C(_06116_),
    .X(_06765_));
 sky130_fd_sc_hd__clkbuf_4 _11721_ (.A(_05996_),
    .X(_06766_));
 sky130_fd_sc_hd__and3_1 _11722_ (.A(\cur_mb_mem[230][5] ),
    .B(_06204_),
    .C(_06766_),
    .X(_06767_));
 sky130_fd_sc_hd__and3_1 _11723_ (.A(\cur_mb_mem[63][5] ),
    .B(_06149_),
    .C(_06198_),
    .X(_06768_));
 sky130_fd_sc_hd__a2111o_2 _11724_ (.A1(\cur_mb_mem[231][5] ),
    .A2(_06180_),
    .B1(_06765_),
    .C1(_06767_),
    .D1(_06768_),
    .X(_06769_));
 sky130_fd_sc_hd__clkbuf_16 _11725_ (.A(_06060_),
    .X(_06770_));
 sky130_fd_sc_hd__and3_1 _11726_ (.A(\cur_mb_mem[227][5] ),
    .B(_06770_),
    .C(_06766_),
    .X(_06771_));
 sky130_fd_sc_hd__clkbuf_16 _11727_ (.A(net237),
    .X(_06772_));
 sky130_fd_sc_hd__and3_1 _11728_ (.A(\cur_mb_mem[224][5] ),
    .B(_06772_),
    .C(_06247_),
    .X(_06773_));
 sky130_fd_sc_hd__clkbuf_16 _11729_ (.A(net256),
    .X(_06774_));
 sky130_fd_sc_hd__clkbuf_4 _11730_ (.A(_05997_),
    .X(_06775_));
 sky130_fd_sc_hd__and3_1 _11731_ (.A(\cur_mb_mem[232][5] ),
    .B(_06774_),
    .C(_06775_),
    .X(_06776_));
 sky130_fd_sc_hd__a2111o_2 _11732_ (.A1(\cur_mb_mem[234][5] ),
    .A2(_06117_),
    .B1(_06771_),
    .C1(_06773_),
    .D1(_06776_),
    .X(_06777_));
 sky130_fd_sc_hd__or4_4 _11733_ (.A(_06757_),
    .B(_06764_),
    .C(_06769_),
    .D(_06777_),
    .X(_06778_));
 sky130_fd_sc_hd__or4_1 _11734_ (.A(_06711_),
    .B(_06730_),
    .C(_06751_),
    .D(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__and3_1 _11735_ (.A(\cur_mb_mem[154][5] ),
    .B(_06442_),
    .C(_06188_),
    .X(_06780_));
 sky130_fd_sc_hd__and3_1 _11736_ (.A(\cur_mb_mem[145][5] ),
    .B(_06188_),
    .C(_06076_),
    .X(_06781_));
 sky130_fd_sc_hd__and3_1 _11737_ (.A(\cur_mb_mem[100][5] ),
    .B(_06744_),
    .C(_06045_),
    .X(_06782_));
 sky130_fd_sc_hd__a2111o_1 _11738_ (.A1(\cur_mb_mem[159][5] ),
    .A2(_06174_),
    .B1(_06780_),
    .C1(_06781_),
    .D1(_06782_),
    .X(_06783_));
 sky130_fd_sc_hd__and3_1 _11739_ (.A(\cur_mb_mem[103][5] ),
    .B(_06027_),
    .C(_06461_),
    .X(_06784_));
 sky130_fd_sc_hd__and3_1 _11740_ (.A(\cur_mb_mem[99][5] ),
    .B(_06313_),
    .C(_06347_),
    .X(_06785_));
 sky130_fd_sc_hd__and3_1 _11741_ (.A(\cur_mb_mem[95][5] ),
    .B(_06120_),
    .C(_06378_),
    .X(_06786_));
 sky130_fd_sc_hd__a2111o_1 _11742_ (.A1(\cur_mb_mem[15][5] ),
    .A2(_06295_),
    .B1(_06784_),
    .C1(_06785_),
    .D1(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__and3_1 _11743_ (.A(\cur_mb_mem[105][5] ),
    .B(_05892_),
    .C(_06267_),
    .X(_06788_));
 sky130_fd_sc_hd__clkbuf_8 _11744_ (.A(_06081_),
    .X(_06789_));
 sky130_fd_sc_hd__and3_1 _11745_ (.A(\cur_mb_mem[207][5] ),
    .B(_06099_),
    .C(_06789_),
    .X(_06790_));
 sky130_fd_sc_hd__and3_1 _11746_ (.A(\cur_mb_mem[96][5] ),
    .B(_06267_),
    .C(net236),
    .X(_06791_));
 sky130_fd_sc_hd__and3_1 _11747_ (.A(\cur_mb_mem[157][5] ),
    .B(_05944_),
    .C(_05977_),
    .X(_06792_));
 sky130_fd_sc_hd__or4_1 _11748_ (.A(_06788_),
    .B(_06790_),
    .C(_06791_),
    .D(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__buf_8 _11749_ (.A(_06130_),
    .X(_06794_));
 sky130_fd_sc_hd__and3_1 _11750_ (.A(\cur_mb_mem[101][5] ),
    .B(_06268_),
    .C(_06794_),
    .X(_06795_));
 sky130_fd_sc_hd__a221o_1 _11751_ (.A1(\cur_mb_mem[153][5] ),
    .A2(_06453_),
    .B1(_06305_),
    .B2(\cur_mb_mem[143][5] ),
    .C1(_06795_),
    .X(_06796_));
 sky130_fd_sc_hd__or4_2 _11752_ (.A(_06783_),
    .B(_06787_),
    .C(_06793_),
    .D(_06796_),
    .X(_06797_));
 sky130_fd_sc_hd__and3_1 _11753_ (.A(\cur_mb_mem[247][5] ),
    .B(_06032_),
    .C(_06461_),
    .X(_06798_));
 sky130_fd_sc_hd__and3_1 _11754_ (.A(\cur_mb_mem[202][5] ),
    .B(_05931_),
    .C(_06324_),
    .X(_06799_));
 sky130_fd_sc_hd__and3_1 _11755_ (.A(\cur_mb_mem[252][5] ),
    .B(_06158_),
    .C(_06718_),
    .X(_06800_));
 sky130_fd_sc_hd__a2111o_1 _11756_ (.A1(\cur_mb_mem[253][5] ),
    .A2(_06034_),
    .B1(_06798_),
    .C1(_06799_),
    .D1(_06800_),
    .X(_06801_));
 sky130_fd_sc_hd__clkbuf_4 _11757_ (.A(_05939_),
    .X(_06802_));
 sky130_fd_sc_hd__and3_1 _11758_ (.A(\cur_mb_mem[212][5] ),
    .B(_06026_),
    .C(_06802_),
    .X(_06803_));
 sky130_fd_sc_hd__and3_1 _11759_ (.A(\cur_mb_mem[220][5] ),
    .B(_06321_),
    .C(_06348_),
    .X(_06804_));
 sky130_fd_sc_hd__and3_1 _11760_ (.A(\cur_mb_mem[104][5] ),
    .B(_06455_),
    .C(_06045_),
    .X(_06805_));
 sky130_fd_sc_hd__a2111o_1 _11761_ (.A1(\cur_mb_mem[250][5] ),
    .A2(_06443_),
    .B1(_06803_),
    .C1(_06804_),
    .D1(_06805_),
    .X(_06806_));
 sky130_fd_sc_hd__and3_1 _11762_ (.A(\cur_mb_mem[245][5] ),
    .B(_06158_),
    .C(_06131_),
    .X(_06807_));
 sky130_fd_sc_hd__and3_1 _11763_ (.A(\cur_mb_mem[193][5] ),
    .B(_06456_),
    .C(_05995_),
    .X(_06808_));
 sky130_fd_sc_hd__buf_6 _11764_ (.A(_06022_),
    .X(_06809_));
 sky130_fd_sc_hd__and3_4 _11765_ (.A(\cur_mb_mem[79][5] ),
    .B(_06466_),
    .C(_06809_),
    .X(_06810_));
 sky130_fd_sc_hd__a2111o_1 _11766_ (.A1(\cur_mb_mem[108][5] ),
    .A2(_06322_),
    .B1(_06807_),
    .C1(_06808_),
    .D1(_06810_),
    .X(_06811_));
 sky130_fd_sc_hd__buf_12 _11767_ (.A(_06130_),
    .X(_06812_));
 sky130_fd_sc_hd__and3_1 _11768_ (.A(\cur_mb_mem[197][5] ),
    .B(_06456_),
    .C(_06812_),
    .X(_06813_));
 sky130_fd_sc_hd__clkbuf_8 _11769_ (.A(_05940_),
    .X(_06814_));
 sky130_fd_sc_hd__buf_12 _11770_ (.A(net239),
    .X(_06815_));
 sky130_fd_sc_hd__and3_1 _11771_ (.A(\cur_mb_mem[208][5] ),
    .B(_06814_),
    .C(_06815_),
    .X(_06816_));
 sky130_fd_sc_hd__and3_1 _11772_ (.A(\cur_mb_mem[205][5] ),
    .B(_06762_),
    .C(_06082_),
    .X(_06817_));
 sky130_fd_sc_hd__a2111o_1 _11773_ (.A1(\cur_mb_mem[111][5] ),
    .A2(_06069_),
    .B1(_06813_),
    .C1(_06816_),
    .D1(_06817_),
    .X(_06818_));
 sky130_fd_sc_hd__or4_4 _11774_ (.A(_06801_),
    .B(_06806_),
    .C(_06811_),
    .D(_06818_),
    .X(_06819_));
 sky130_fd_sc_hd__a32o_1 _11775_ (.A1(\cur_mb_mem[13][5] ),
    .A2(_06112_),
    .A3(_05946_),
    .B1(_06284_),
    .B2(\cur_mb_mem[162][5] ),
    .X(_06820_));
 sky130_fd_sc_hd__a32o_1 _11776_ (.A1(\cur_mb_mem[167][5] ),
    .A2(_06137_),
    .A3(_06097_),
    .B1(_06236_),
    .B2(\cur_mb_mem[21][5] ),
    .X(_06821_));
 sky130_fd_sc_hd__or2_1 _11777_ (.A(_06820_),
    .B(_06821_),
    .X(_06822_));
 sky130_fd_sc_hd__a32o_2 _11778_ (.A1(\cur_mb_mem[213][5] ),
    .A2(_05941_),
    .A3(_06132_),
    .B1(_06193_),
    .B2(\cur_mb_mem[166][5] ),
    .X(_06823_));
 sky130_fd_sc_hd__a32o_2 _11779_ (.A1(\cur_mb_mem[20][5] ),
    .A2(_06134_),
    .A3(_05975_),
    .B1(_06301_),
    .B2(\cur_mb_mem[11][5] ),
    .X(_06824_));
 sky130_fd_sc_hd__clkbuf_8 _11780_ (.A(_05921_),
    .X(_06825_));
 sky130_fd_sc_hd__and3_1 _11781_ (.A(\cur_mb_mem[165][5] ),
    .B(_06825_),
    .C(_06812_),
    .X(_06826_));
 sky130_fd_sc_hd__and3_1 _11782_ (.A(\cur_mb_mem[6][5] ),
    .B(_06707_),
    .C(_06199_),
    .X(_06827_));
 sky130_fd_sc_hd__and3_1 _11783_ (.A(\cur_mb_mem[160][5] ),
    .B(_06192_),
    .C(_06748_),
    .X(_06828_));
 sky130_fd_sc_hd__a2111o_1 _11784_ (.A1(\cur_mb_mem[73][5] ),
    .A2(_06328_),
    .B1(_06826_),
    .C1(_06827_),
    .D1(_06828_),
    .X(_06829_));
 sky130_fd_sc_hd__buf_6 _11785_ (.A(_06018_),
    .X(_06830_));
 sky130_fd_sc_hd__and3_1 _11786_ (.A(\cur_mb_mem[186][5] ),
    .B(_05957_),
    .C(_06830_),
    .X(_06831_));
 sky130_fd_sc_hd__buf_12 _11787_ (.A(net2007),
    .X(_06832_));
 sky130_fd_sc_hd__and3_1 _11788_ (.A(\cur_mb_mem[184][5] ),
    .B(_06832_),
    .C(_06830_),
    .X(_06833_));
 sky130_fd_sc_hd__buf_8 _11789_ (.A(_05892_),
    .X(_06834_));
 sky130_fd_sc_hd__and3_1 _11790_ (.A(\cur_mb_mem[185][5] ),
    .B(_06834_),
    .C(_06216_),
    .X(_06835_));
 sky130_fd_sc_hd__a2111o_1 _11791_ (.A1(\cur_mb_mem[74][5] ),
    .A2(_06417_),
    .B1(_06831_),
    .C1(_06833_),
    .D1(_06835_),
    .X(_06836_));
 sky130_fd_sc_hd__or4_1 _11792_ (.A(_06823_),
    .B(_06824_),
    .C(_06829_),
    .D(_06836_),
    .X(_06837_));
 sky130_fd_sc_hd__or4_1 _11793_ (.A(_06797_),
    .B(_06819_),
    .C(_06822_),
    .D(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__and3_1 _11794_ (.A(\cur_mb_mem[183][5] ),
    .B(_06013_),
    .C(_06461_),
    .X(_06839_));
 sky130_fd_sc_hd__and3_1 _11795_ (.A(\cur_mb_mem[131][5] ),
    .B(_06347_),
    .C(_05933_),
    .X(_06840_));
 sky130_fd_sc_hd__buf_12 _11796_ (.A(net231),
    .X(_06841_));
 sky130_fd_sc_hd__clkbuf_8 _11797_ (.A(net248),
    .X(_06842_));
 sky130_fd_sc_hd__and3_1 _11798_ (.A(\cur_mb_mem[129][5] ),
    .B(_06841_),
    .C(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__a2111o_1 _11799_ (.A1(\cur_mb_mem[128][5] ),
    .A2(_06075_),
    .B1(_06839_),
    .C1(_06840_),
    .D1(_06843_),
    .X(_06844_));
 sky130_fd_sc_hd__and3_1 _11800_ (.A(\cur_mb_mem[182][5] ),
    .B(_06210_),
    .C(_06013_),
    .X(_06845_));
 sky130_fd_sc_hd__and3_1 _11801_ (.A(\cur_mb_mem[57][5] ),
    .B(_06170_),
    .C(_06038_),
    .X(_06846_));
 sky130_fd_sc_hd__and3_2 _11802_ (.A(\cur_mb_mem[107][5] ),
    .B(_06474_),
    .C(_05984_),
    .X(_06847_));
 sky130_fd_sc_hd__a2111o_1 _11803_ (.A1(\cur_mb_mem[135][5] ),
    .A2(_06462_),
    .B1(_06845_),
    .C1(_06846_),
    .D1(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__clkbuf_8 _11804_ (.A(_05055_),
    .X(_06849_));
 sky130_fd_sc_hd__and3_1 _11805_ (.A(\cur_mb_mem[60][5] ),
    .B(_06849_),
    .C(_05901_),
    .X(_06850_));
 sky130_fd_sc_hd__clkbuf_16 _11806_ (.A(_06095_),
    .X(_06851_));
 sky130_fd_sc_hd__and3_1 _11807_ (.A(\cur_mb_mem[55][5] ),
    .B(_06849_),
    .C(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__and3_1 _11808_ (.A(\cur_mb_mem[178][5] ),
    .B(_06079_),
    .C(_06018_),
    .X(_06853_));
 sky130_fd_sc_hd__and3_1 _11809_ (.A(\cur_mb_mem[177][5] ),
    .B(_06013_),
    .C(net230),
    .X(_06854_));
 sky130_fd_sc_hd__or4_1 _11810_ (.A(_06850_),
    .B(_06852_),
    .C(_06853_),
    .D(_06854_),
    .X(_06855_));
 sky130_fd_sc_hd__clkbuf_8 _11811_ (.A(_05055_),
    .X(_06856_));
 sky130_fd_sc_hd__and3_1 _11812_ (.A(\cur_mb_mem[49][5] ),
    .B(_06856_),
    .C(_06353_),
    .X(_06857_));
 sky130_fd_sc_hd__and3_1 _11813_ (.A(\cur_mb_mem[36][5] ),
    .B(_06232_),
    .C(_06343_),
    .X(_06858_));
 sky130_fd_sc_hd__buf_8 _11814_ (.A(net248),
    .X(_06859_));
 sky130_fd_sc_hd__and3_1 _11815_ (.A(\cur_mb_mem[134][5] ),
    .B(_06191_),
    .C(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__a2111o_1 _11816_ (.A1(\cur_mb_mem[50][5] ),
    .A2(_06172_),
    .B1(_06857_),
    .C1(_06858_),
    .D1(_06860_),
    .X(_06861_));
 sky130_fd_sc_hd__or4_4 _11817_ (.A(_06844_),
    .B(_06848_),
    .C(_06855_),
    .D(_06861_),
    .X(_06862_));
 sky130_fd_sc_hd__and3_1 _11818_ (.A(\cur_mb_mem[31][5] ),
    .B(_06068_),
    .C(_06403_),
    .X(_06863_));
 sky130_fd_sc_hd__and3_2 _11819_ (.A(\cur_mb_mem[223][5] ),
    .B(_06120_),
    .C(_06348_),
    .X(_06864_));
 sky130_fd_sc_hd__and3_1 _11820_ (.A(\cur_mb_mem[163][5] ),
    .B(_06289_),
    .C(_06825_),
    .X(_06865_));
 sky130_fd_sc_hd__a2111o_1 _11821_ (.A1(\cur_mb_mem[47][5] ),
    .A2(_06259_),
    .B1(_06863_),
    .C1(_06864_),
    .D1(_06865_),
    .X(_06866_));
 sky130_fd_sc_hd__and3_4 _11822_ (.A(\cur_mb_mem[198][5] ),
    .B(_06210_),
    .C(_06324_),
    .X(_06867_));
 sky130_fd_sc_hd__and3_1 _11823_ (.A(\cur_mb_mem[102][5] ),
    .B(_06313_),
    .C(_06210_),
    .X(_06868_));
 sky130_fd_sc_hd__and3_1 _11824_ (.A(\cur_mb_mem[106][5] ),
    .B(_05957_),
    .C(_05984_),
    .X(_06869_));
 sky130_fd_sc_hd__a2111o_1 _11825_ (.A1(\cur_mb_mem[98][5] ),
    .A2(_06330_),
    .B1(_06867_),
    .C1(_06868_),
    .D1(_06869_),
    .X(_06870_));
 sky130_fd_sc_hd__and3_1 _11826_ (.A(\cur_mb_mem[175][5] ),
    .B(_06068_),
    .C(_06333_),
    .X(_06871_));
 sky130_fd_sc_hd__and3_1 _11827_ (.A(\cur_mb_mem[161][5] ),
    .B(_05995_),
    .C(_06825_),
    .X(_06872_));
 sky130_fd_sc_hd__and3_1 _11828_ (.A(\cur_mb_mem[180][5] ),
    .B(_06232_),
    .C(_06760_),
    .X(_06873_));
 sky130_fd_sc_hd__a2111o_1 _11829_ (.A1(\cur_mb_mem[97][5] ),
    .A2(_06077_),
    .B1(_06871_),
    .C1(_06872_),
    .D1(_06873_),
    .X(_06874_));
 sky130_fd_sc_hd__and3_1 _11830_ (.A(\cur_mb_mem[109][5] ),
    .B(_05984_),
    .C(_06490_),
    .X(_06875_));
 sky130_fd_sc_hd__and3_1 _11831_ (.A(\cur_mb_mem[148][5] ),
    .B(_06232_),
    .C(_06401_),
    .X(_06876_));
 sky130_fd_sc_hd__clkbuf_16 _11832_ (.A(_06018_),
    .X(_06877_));
 sky130_fd_sc_hd__and3_1 _11833_ (.A(\cur_mb_mem[181][5] ),
    .B(_06877_),
    .C(_06794_),
    .X(_06878_));
 sky130_fd_sc_hd__a2111o_1 _11834_ (.A1(\cur_mb_mem[110][5] ),
    .A2(_06047_),
    .B1(_06875_),
    .C1(_06876_),
    .D1(_06878_),
    .X(_06879_));
 sky130_fd_sc_hd__or4_1 _11835_ (.A(_06866_),
    .B(_06870_),
    .C(_06874_),
    .D(_06879_),
    .X(_06880_));
 sky130_fd_sc_hd__and3_1 _11836_ (.A(\cur_mb_mem[48][5] ),
    .B(_06170_),
    .C(_06009_),
    .X(_06881_));
 sky130_fd_sc_hd__and3_1 _11837_ (.A(\cur_mb_mem[71][5] ),
    .B(_06121_),
    .C(_06179_),
    .X(_06882_));
 sky130_fd_sc_hd__and3_1 _11838_ (.A(\cur_mb_mem[64][5] ),
    .B(_06809_),
    .C(_05970_),
    .X(_06883_));
 sky130_fd_sc_hd__a2111o_1 _11839_ (.A1(\cur_mb_mem[65][5] ),
    .A2(_06483_),
    .B1(_06881_),
    .C1(_06882_),
    .D1(_06883_),
    .X(_06884_));
 sky130_fd_sc_hd__and3_1 _11840_ (.A(\cur_mb_mem[62][5] ),
    .B(_06170_),
    .C(_06046_),
    .X(_06885_));
 sky130_fd_sc_hd__and3_1 _11841_ (.A(\cur_mb_mem[58][5] ),
    .B(_06350_),
    .C(_06115_),
    .X(_06886_));
 sky130_fd_sc_hd__and3_1 _11842_ (.A(\cur_mb_mem[141][5] ),
    .B(_06762_),
    .C(_06842_),
    .X(_06887_));
 sky130_fd_sc_hd__a2111o_1 _11843_ (.A1(\cur_mb_mem[140][5] ),
    .A2(_06423_),
    .B1(_06885_),
    .C1(_06886_),
    .D1(_06887_),
    .X(_06888_));
 sky130_fd_sc_hd__and3_1 _11844_ (.A(\cur_mb_mem[44][5] ),
    .B(_06422_),
    .C(_06395_),
    .X(_06889_));
 sky130_fd_sc_hd__and3_1 _11845_ (.A(\cur_mb_mem[176][5] ),
    .B(_06019_),
    .C(_06815_),
    .X(_06890_));
 sky130_fd_sc_hd__and3_1 _11846_ (.A(\cur_mb_mem[56][5] ),
    .B(_06240_),
    .C(_05982_),
    .X(_06891_));
 sky130_fd_sc_hd__a2111o_2 _11847_ (.A1(\cur_mb_mem[61][5] ),
    .A2(_06359_),
    .B1(_06889_),
    .C1(_06890_),
    .D1(_06891_),
    .X(_06892_));
 sky130_fd_sc_hd__and3_1 _11848_ (.A(\cur_mb_mem[86][5] ),
    .B(_05914_),
    .C(_06204_),
    .X(_06893_));
 sky130_fd_sc_hd__and3_1 _11849_ (.A(\cur_mb_mem[93][5] ),
    .B(_06230_),
    .C(_06762_),
    .X(_06894_));
 sky130_fd_sc_hd__buf_8 _11850_ (.A(net253),
    .X(_06895_));
 sky130_fd_sc_hd__buf_8 _11851_ (.A(_06095_),
    .X(_06896_));
 sky130_fd_sc_hd__and3_1 _11852_ (.A(\cur_mb_mem[87][5] ),
    .B(_06895_),
    .C(_06896_),
    .X(_06897_));
 sky130_fd_sc_hd__a2111o_1 _11853_ (.A1(\cur_mb_mem[80][5] ),
    .A2(_06010_),
    .B1(_06893_),
    .C1(_06894_),
    .D1(_06897_),
    .X(_06898_));
 sky130_fd_sc_hd__or4_4 _11854_ (.A(_06884_),
    .B(_06888_),
    .C(_06892_),
    .D(_06898_),
    .X(_06899_));
 sky130_fd_sc_hd__and3_1 _11855_ (.A(\cur_mb_mem[235][5] ),
    .B(_06312_),
    .C(_06116_),
    .X(_06900_));
 sky130_fd_sc_hd__and3_1 _11856_ (.A(\cur_mb_mem[240][5] ),
    .B(_06165_),
    .C(_05970_),
    .X(_06901_));
 sky130_fd_sc_hd__clkbuf_8 _11857_ (.A(_04429_),
    .X(_06902_));
 sky130_fd_sc_hd__buf_8 _11858_ (.A(_05892_),
    .X(_06903_));
 sky130_fd_sc_hd__and3_1 _11859_ (.A(\cur_mb_mem[249][5] ),
    .B(_06902_),
    .C(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__a2111o_1 _11860_ (.A1(\cur_mb_mem[248][5] ),
    .A2(_06411_),
    .B1(_06900_),
    .C1(_06901_),
    .D1(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__and3_1 _11861_ (.A(\cur_mb_mem[251][5] ),
    .B(_06165_),
    .C(_06312_),
    .X(_06906_));
 sky130_fd_sc_hd__and3_1 _11862_ (.A(\cur_mb_mem[59][5] ),
    .B(_06240_),
    .C(_06474_),
    .X(_06907_));
 sky130_fd_sc_hd__clkbuf_16 _11863_ (.A(_06078_),
    .X(_06908_));
 sky130_fd_sc_hd__and3_1 _11864_ (.A(\cur_mb_mem[242][5] ),
    .B(_06902_),
    .C(_06908_),
    .X(_06909_));
 sky130_fd_sc_hd__a2111o_1 _11865_ (.A1(\cur_mb_mem[246][5] ),
    .A2(_06160_),
    .B1(_06906_),
    .C1(_06907_),
    .D1(_06909_),
    .X(_06910_));
 sky130_fd_sc_hd__and3_1 _11866_ (.A(\cur_mb_mem[228][5] ),
    .B(_06232_),
    .C(_06255_),
    .X(_06911_));
 sky130_fd_sc_hd__buf_12 _11867_ (.A(net230),
    .X(_06912_));
 sky130_fd_sc_hd__and3_1 _11868_ (.A(\cur_mb_mem[225][5] ),
    .B(_06912_),
    .C(_06766_),
    .X(_06913_));
 sky130_fd_sc_hd__and3_1 _11869_ (.A(\cur_mb_mem[254][5] ),
    .B(_06902_),
    .C(_06000_),
    .X(_06914_));
 sky130_fd_sc_hd__a2111o_1 _11870_ (.A1(\cur_mb_mem[255][5] ),
    .A2(_06304_),
    .B1(_06911_),
    .C1(_06913_),
    .D1(_06914_),
    .X(_06915_));
 sky130_fd_sc_hd__clkbuf_8 _11871_ (.A(_04429_),
    .X(_06916_));
 sky130_fd_sc_hd__and3_1 _11872_ (.A(\cur_mb_mem[243][5] ),
    .B(_06916_),
    .C(_06770_),
    .X(_06917_));
 sky130_fd_sc_hd__buf_4 _11873_ (.A(_05997_),
    .X(_06918_));
 sky130_fd_sc_hd__and3_1 _11874_ (.A(\cur_mb_mem[226][5] ),
    .B(_06908_),
    .C(_06918_),
    .X(_06919_));
 sky130_fd_sc_hd__clkbuf_16 _11875_ (.A(_05901_),
    .X(_06920_));
 sky130_fd_sc_hd__and3_1 _11876_ (.A(\cur_mb_mem[236][5] ),
    .B(_06920_),
    .C(_06775_),
    .X(_06921_));
 sky130_fd_sc_hd__a2111o_1 _11877_ (.A1(\cur_mb_mem[127][5] ),
    .A2(_06101_),
    .B1(_06917_),
    .C1(_06919_),
    .D1(_06921_),
    .X(_06922_));
 sky130_fd_sc_hd__or4_4 _11878_ (.A(_06905_),
    .B(_06910_),
    .C(_06915_),
    .D(_06922_),
    .X(_06923_));
 sky130_fd_sc_hd__or4_1 _11879_ (.A(_06862_),
    .B(_06880_),
    .C(_06899_),
    .D(_06923_),
    .X(_06924_));
 sky130_fd_sc_hd__and3_1 _11880_ (.A(\cur_mb_mem[94][5] ),
    .B(_06008_),
    .C(_06435_),
    .X(_06925_));
 sky130_fd_sc_hd__and3_1 _11881_ (.A(\cur_mb_mem[68][5] ),
    .B(_06166_),
    .C(_06233_),
    .X(_06926_));
 sky130_fd_sc_hd__clkbuf_8 _11882_ (.A(net253),
    .X(_06927_));
 sky130_fd_sc_hd__and3_1 _11883_ (.A(\cur_mb_mem[91][5] ),
    .B(_06400_),
    .C(_06927_),
    .X(_06928_));
 sky130_fd_sc_hd__a2111o_1 _11884_ (.A1(\cur_mb_mem[136][5] ),
    .A2(_06292_),
    .B1(_06925_),
    .C1(_06926_),
    .D1(_06928_),
    .X(_06929_));
 sky130_fd_sc_hd__and3_1 _11885_ (.A(\cur_mb_mem[69][5] ),
    .B(_06121_),
    .C(_06220_),
    .X(_06930_));
 sky130_fd_sc_hd__clkbuf_16 _11886_ (.A(_05913_),
    .X(_06931_));
 sky130_fd_sc_hd__and3_1 _11887_ (.A(\cur_mb_mem[90][5] ),
    .B(_06115_),
    .C(_06931_),
    .X(_06932_));
 sky130_fd_sc_hd__and3_4 _11888_ (.A(\cur_mb_mem[219][5] ),
    .B(_06387_),
    .C(_06150_),
    .X(_06933_));
 sky130_fd_sc_hd__a2111o_1 _11889_ (.A1(\cur_mb_mem[40][5] ),
    .A2(_06485_),
    .B1(_06930_),
    .C1(_06932_),
    .D1(_06933_),
    .X(_06934_));
 sky130_fd_sc_hd__and3_1 _11890_ (.A(\cur_mb_mem[46][5] ),
    .B(_06343_),
    .C(_06435_),
    .X(_06935_));
 sky130_fd_sc_hd__and3_1 _11891_ (.A(\cur_mb_mem[83][5] ),
    .B(_05914_),
    .C(_06289_),
    .X(_06936_));
 sky130_fd_sc_hd__buf_8 _11892_ (.A(_05901_),
    .X(_06937_));
 sky130_fd_sc_hd__and3_1 _11893_ (.A(\cur_mb_mem[92][5] ),
    .B(_06937_),
    .C(_06927_),
    .X(_06938_));
 sky130_fd_sc_hd__a2111o_1 _11894_ (.A1(\cur_mb_mem[70][5] ),
    .A2(_06144_),
    .B1(_06935_),
    .C1(_06936_),
    .D1(_06938_),
    .X(_06939_));
 sky130_fd_sc_hd__and3_1 _11895_ (.A(\cur_mb_mem[81][5] ),
    .B(_06230_),
    .C(_06841_),
    .X(_06940_));
 sky130_fd_sc_hd__and3_1 _11896_ (.A(\cur_mb_mem[82][5] ),
    .B(_06908_),
    .C(_06927_),
    .X(_06941_));
 sky130_fd_sc_hd__clkbuf_16 _11897_ (.A(_05917_),
    .X(_06942_));
 sky130_fd_sc_hd__and3_1 _11898_ (.A(\cur_mb_mem[139][5] ),
    .B(_06942_),
    .C(_06859_),
    .X(_06943_));
 sky130_fd_sc_hd__a2111o_1 _11899_ (.A1(\cur_mb_mem[45][5] ),
    .A2(_06491_),
    .B1(_06940_),
    .C1(_06941_),
    .D1(_06943_),
    .X(_06944_));
 sky130_fd_sc_hd__or4_4 _11900_ (.A(_06929_),
    .B(_06934_),
    .C(_06939_),
    .D(_06944_),
    .X(_06945_));
 sky130_fd_sc_hd__and3_1 _11901_ (.A(\cur_mb_mem[130][5] ),
    .B(_06341_),
    .C(_06382_),
    .X(_06946_));
 sky130_fd_sc_hd__and3_1 _11902_ (.A(\cur_mb_mem[52][5] ),
    .B(_06856_),
    .C(_06166_),
    .X(_06947_));
 sky130_fd_sc_hd__and3_1 _11903_ (.A(\cur_mb_mem[54][5] ),
    .B(_06198_),
    .C(_06199_),
    .X(_06948_));
 sky130_fd_sc_hd__a2111o_4 _11904_ (.A1(\cur_mb_mem[53][5] ),
    .A2(_06221_),
    .B1(_06946_),
    .C1(_06947_),
    .D1(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__and3_1 _11905_ (.A(\cur_mb_mem[51][5] ),
    .B(_06350_),
    .C(_06355_),
    .X(_06950_));
 sky130_fd_sc_hd__and3_1 _11906_ (.A(\cur_mb_mem[229][5] ),
    .B(_06147_),
    .C(_06255_),
    .X(_06951_));
 sky130_fd_sc_hd__buf_6 _11907_ (.A(net2004),
    .X(_06952_));
 sky130_fd_sc_hd__and3_1 _11908_ (.A(\cur_mb_mem[39][5] ),
    .B(_06952_),
    .C(_06708_),
    .X(_06953_));
 sky130_fd_sc_hd__a2111o_1 _11909_ (.A1(\cur_mb_mem[38][5] ),
    .A2(_06396_),
    .B1(_06950_),
    .C1(_06951_),
    .D1(_06953_),
    .X(_06954_));
 sky130_fd_sc_hd__and3_1 _11910_ (.A(\cur_mb_mem[191][5] ),
    .B(_06466_),
    .C(_06019_),
    .X(_06955_));
 sky130_fd_sc_hd__and3_1 _11911_ (.A(\cur_mb_mem[216][5] ),
    .B(_06478_),
    .C(_06814_),
    .X(_06956_));
 sky130_fd_sc_hd__and3_1 _11912_ (.A(\cur_mb_mem[37][5] ),
    .B(_06087_),
    .C(_06794_),
    .X(_06957_));
 sky130_fd_sc_hd__a2111o_1 _11913_ (.A1(\cur_mb_mem[239][5] ),
    .A2(_06125_),
    .B1(_06955_),
    .C1(_06956_),
    .D1(_06957_),
    .X(_06958_));
 sky130_fd_sc_hd__and3_2 _11914_ (.A(\cur_mb_mem[241][5] ),
    .B(_06916_),
    .C(_06912_),
    .X(_06959_));
 sky130_fd_sc_hd__clkbuf_16 _11915_ (.A(_05904_),
    .X(_06960_));
 sky130_fd_sc_hd__and3_1 _11916_ (.A(\cur_mb_mem[218][5] ),
    .B(_06960_),
    .C(_06150_),
    .X(_06961_));
 sky130_fd_sc_hd__and3_1 _11917_ (.A(\cur_mb_mem[210][5] ),
    .B(_06380_),
    .C(_05947_),
    .X(_06962_));
 sky130_fd_sc_hd__a2111o_4 _11918_ (.A1(\cur_mb_mem[209][5] ),
    .A2(_06271_),
    .B1(_06959_),
    .C1(_06961_),
    .D1(_06962_),
    .X(_06963_));
 sky130_fd_sc_hd__or4_4 _11919_ (.A(_06949_),
    .B(_06954_),
    .C(_06958_),
    .D(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__and3_1 _11920_ (.A(\cur_mb_mem[214][5] ),
    .B(_06140_),
    .C(_06270_),
    .X(_06965_));
 sky130_fd_sc_hd__and3_1 _11921_ (.A(\cur_mb_mem[170][5] ),
    .B(_05957_),
    .C(_06825_),
    .X(_06966_));
 sky130_fd_sc_hd__buf_8 _11922_ (.A(_06081_),
    .X(_06967_));
 sky130_fd_sc_hd__and3_1 _11923_ (.A(\cur_mb_mem[199][5] ),
    .B(_06967_),
    .C(_06896_),
    .X(_06968_));
 sky130_fd_sc_hd__a2111o_4 _11924_ (.A1(\cur_mb_mem[200][5] ),
    .A2(_06457_),
    .B1(_06965_),
    .C1(_06966_),
    .D1(_06968_),
    .X(_06969_));
 sky130_fd_sc_hd__and3_1 _11925_ (.A(\cur_mb_mem[169][5] ),
    .B(_05892_),
    .C(_05921_),
    .X(_06970_));
 sky130_fd_sc_hd__and3_1 _11926_ (.A(\cur_mb_mem[222][5] ),
    .B(_05940_),
    .C(_05953_),
    .X(_06971_));
 sky130_fd_sc_hd__and3_1 _11927_ (.A(\cur_mb_mem[221][5] ),
    .B(_06033_),
    .C(_05940_),
    .X(_06972_));
 sky130_fd_sc_hd__and3_2 _11928_ (.A(\cur_mb_mem[32][5] ),
    .B(_06005_),
    .C(_06074_),
    .X(_06973_));
 sky130_fd_sc_hd__or4_4 _11929_ (.A(_06970_),
    .B(_06971_),
    .C(_06972_),
    .D(_06973_),
    .X(_06974_));
 sky130_fd_sc_hd__and3_1 _11930_ (.A(\cur_mb_mem[88][5] ),
    .B(_06478_),
    .C(_05914_),
    .X(_06975_));
 sky130_fd_sc_hd__and3_1 _11931_ (.A(\cur_mb_mem[137][5] ),
    .B(_06903_),
    .C(_06842_),
    .X(_06976_));
 sky130_fd_sc_hd__and3_1 _11932_ (.A(\cur_mb_mem[33][5] ),
    .B(_06087_),
    .C(_06251_),
    .X(_06977_));
 sky130_fd_sc_hd__a2111o_1 _11933_ (.A1(\cur_mb_mem[215][5] ),
    .A2(_06447_),
    .B1(_06975_),
    .C1(_06976_),
    .D1(_06977_),
    .X(_06978_));
 sky130_fd_sc_hd__and3_1 _11934_ (.A(\cur_mb_mem[89][5] ),
    .B(_06903_),
    .C(_06927_),
    .X(_06979_));
 sky130_fd_sc_hd__clkbuf_16 _11935_ (.A(_06061_),
    .X(_06980_));
 sky130_fd_sc_hd__and3_1 _11936_ (.A(\cur_mb_mem[35][5] ),
    .B(_06980_),
    .C(_06087_),
    .X(_06981_));
 sky130_fd_sc_hd__and3_1 _11937_ (.A(\cur_mb_mem[138][5] ),
    .B(_05905_),
    .C(_05935_),
    .X(_06982_));
 sky130_fd_sc_hd__a2111o_1 _11938_ (.A1(\cur_mb_mem[34][5] ),
    .A2(_06393_),
    .B1(_06979_),
    .C1(_06981_),
    .D1(_06982_),
    .X(_06983_));
 sky130_fd_sc_hd__or4_1 _11939_ (.A(_06969_),
    .B(_06974_),
    .C(_06978_),
    .D(_06983_),
    .X(_06984_));
 sky130_fd_sc_hd__and3_1 _11940_ (.A(\cur_mb_mem[168][5] ),
    .B(_05895_),
    .C(_06333_),
    .X(_06985_));
 sky130_fd_sc_hd__clkbuf_4 _11941_ (.A(_06081_),
    .X(_06986_));
 sky130_fd_sc_hd__and3_1 _11942_ (.A(\cur_mb_mem[194][5] ),
    .B(_06079_),
    .C(_06986_),
    .X(_06987_));
 sky130_fd_sc_hd__and3_1 _11943_ (.A(\cur_mb_mem[204][5] ),
    .B(_06321_),
    .C(_06986_),
    .X(_06988_));
 sky130_fd_sc_hd__and3_1 _11944_ (.A(\cur_mb_mem[211][5] ),
    .B(_06347_),
    .C(_06348_),
    .X(_06989_));
 sky130_fd_sc_hd__or4_1 _11945_ (.A(_06985_),
    .B(_06987_),
    .C(_06988_),
    .D(_06989_),
    .X(_06990_));
 sky130_fd_sc_hd__and3_1 _11946_ (.A(\cur_mb_mem[195][5] ),
    .B(_06061_),
    .C(_06986_),
    .X(_06991_));
 sky130_fd_sc_hd__and3_1 _11947_ (.A(\cur_mb_mem[142][5] ),
    .B(_06366_),
    .C(_05933_),
    .X(_06992_));
 sky130_fd_sc_hd__and3_1 _11948_ (.A(\cur_mb_mem[217][5] ),
    .B(_05909_),
    .C(_06802_),
    .X(_06993_));
 sky130_fd_sc_hd__and3_1 _11949_ (.A(\cur_mb_mem[201][5] ),
    .B(_06038_),
    .C(_06324_),
    .X(_06994_));
 sky130_fd_sc_hd__or4_1 _11950_ (.A(_06991_),
    .B(_06992_),
    .C(_06993_),
    .D(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__and3_1 _11951_ (.A(\cur_mb_mem[206][5] ),
    .B(_06000_),
    .C(_06082_),
    .X(_06996_));
 sky130_fd_sc_hd__clkbuf_8 _11952_ (.A(_06789_),
    .X(_06997_));
 sky130_fd_sc_hd__and3_1 _11953_ (.A(\cur_mb_mem[192][5] ),
    .B(_06997_),
    .C(_06748_),
    .X(_06998_));
 sky130_fd_sc_hd__and3_2 _11954_ (.A(\cur_mb_mem[237][5] ),
    .B(_06246_),
    .C(_06775_),
    .X(_06999_));
 sky130_fd_sc_hd__a2111o_1 _11955_ (.A1(\cur_mb_mem[244][5] ),
    .A2(_06167_),
    .B1(_06996_),
    .C1(_06998_),
    .D1(_06999_),
    .X(_07000_));
 sky130_fd_sc_hd__buf_8 _11956_ (.A(_05921_),
    .X(_07001_));
 sky130_fd_sc_hd__and3_1 _11957_ (.A(\cur_mb_mem[171][5] ),
    .B(_06942_),
    .C(_07001_),
    .X(_07002_));
 sky130_fd_sc_hd__and3_1 _11958_ (.A(\cur_mb_mem[196][5] ),
    .B(_06215_),
    .C(_06091_),
    .X(_07003_));
 sky130_fd_sc_hd__and3_1 _11959_ (.A(\cur_mb_mem[238][5] ),
    .B(_05954_),
    .C(_06065_),
    .X(_07004_));
 sky130_fd_sc_hd__a2111o_1 _11960_ (.A1(\cur_mb_mem[203][5] ),
    .A2(_06325_),
    .B1(_07002_),
    .C1(_07003_),
    .D1(_07004_),
    .X(_07005_));
 sky130_fd_sc_hd__or4_4 _11961_ (.A(_06990_),
    .B(_06995_),
    .C(_07000_),
    .D(_07005_),
    .X(_07006_));
 sky130_fd_sc_hd__or4_1 _11962_ (.A(_06945_),
    .B(_06964_),
    .C(_06984_),
    .D(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__or4_4 _11963_ (.A(_06779_),
    .B(_06838_),
    .C(_06924_),
    .D(_07007_),
    .X(_07008_));
 sky130_fd_sc_hd__o22ai_4 _11964_ (.A1(\cur_mb_mem[0][5] ),
    .A2(_05908_),
    .B1(_06692_),
    .B2(_07008_),
    .Y(_07009_));
 sky130_fd_sc_hd__nor2_1 _11965_ (.A(net102),
    .B(_07009_),
    .Y(_07010_));
 sky130_fd_sc_hd__a22o_1 _11966_ (.A1(\cur_mb_mem[223][1] ),
    .A2(_06151_),
    .B1(_06297_),
    .B2(\cur_mb_mem[95][1] ),
    .X(_07011_));
 sky130_fd_sc_hd__a32o_2 _11967_ (.A1(\cur_mb_mem[99][1] ),
    .A2(_06299_),
    .A3(_06064_),
    .B1(_06443_),
    .B2(\cur_mb_mem[250][1] ),
    .X(_07012_));
 sky130_fd_sc_hd__a32o_4 _11968_ (.A1(\cur_mb_mem[154][1] ),
    .A2(_05959_),
    .A3(_05979_),
    .B1(_06453_),
    .B2(\cur_mb_mem[153][1] ),
    .X(_07013_));
 sky130_fd_sc_hd__a221o_1 _11969_ (.A1(\cur_mb_mem[28][1] ),
    .A2(_06017_),
    .B1(_06411_),
    .B2(\cur_mb_mem[248][1] ),
    .C1(_07013_),
    .X(_07014_));
 sky130_fd_sc_hd__a211o_1 _11970_ (.A1(\cur_mb_mem[31][1] ),
    .A2(_06178_),
    .B1(_07012_),
    .C1(_07014_),
    .X(_07015_));
 sky130_fd_sc_hd__a32o_1 _11971_ (.A1(\cur_mb_mem[168][1] ),
    .A2(_05896_),
    .A3(_06426_),
    .B1(_06480_),
    .B2(\cur_mb_mem[190][1] ),
    .X(_07016_));
 sky130_fd_sc_hd__a32o_1 _11972_ (.A1(\cur_mb_mem[170][1] ),
    .A2(_05958_),
    .A3(_05923_),
    .B1(_06239_),
    .B2(\cur_mb_mem[116][1] ),
    .X(_07017_));
 sky130_fd_sc_hd__a221o_1 _11973_ (.A1(\cur_mb_mem[98][1] ),
    .A2(_06330_),
    .B1(_06457_),
    .B2(\cur_mb_mem[200][1] ),
    .C1(_07017_),
    .X(_07018_));
 sky130_fd_sc_hd__a22o_1 _11974_ (.A1(\cur_mb_mem[216][1] ),
    .A2(_06317_),
    .B1(_06010_),
    .B2(\cur_mb_mem[80][1] ),
    .X(_07019_));
 sky130_fd_sc_hd__a22o_2 _11975_ (.A1(\cur_mb_mem[24][1] ),
    .A2(_06285_),
    .B1(_06002_),
    .B2(\cur_mb_mem[30][1] ),
    .X(_07020_));
 sky130_fd_sc_hd__buf_8 _11976_ (.A(_06731_),
    .X(_07021_));
 sky130_fd_sc_hd__and3_1 _11977_ (.A(\cur_mb_mem[113][1] ),
    .B(_07021_),
    .C(_05993_),
    .X(_07022_));
 sky130_fd_sc_hd__a31o_1 _11978_ (.A1(\cur_mb_mem[249][1] ),
    .A2(_04430_),
    .A3(_05910_),
    .B1(_07022_),
    .X(_07023_));
 sky130_fd_sc_hd__a32o_1 _11979_ (.A1(\cur_mb_mem[254][1] ),
    .A2(_04430_),
    .A3(_05954_),
    .B1(_06277_),
    .B2(\cur_mb_mem[8][1] ),
    .X(_07024_));
 sky130_fd_sc_hd__a22o_1 _11980_ (.A1(\cur_mb_mem[246][1] ),
    .A2(_06160_),
    .B1(_06047_),
    .B2(\cur_mb_mem[110][1] ),
    .X(_07025_));
 sky130_fd_sc_hd__or4_1 _11981_ (.A(_07020_),
    .B(_07023_),
    .C(_07024_),
    .D(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__or4_2 _11982_ (.A(_07016_),
    .B(_07018_),
    .C(_07019_),
    .D(_07026_),
    .X(_07027_));
 sky130_fd_sc_hd__a2111o_4 _11983_ (.A1(\cur_mb_mem[159][1] ),
    .A2(_06174_),
    .B1(_07011_),
    .C1(_07015_),
    .D1(_07027_),
    .X(_07028_));
 sky130_fd_sc_hd__and3_2 _11984_ (.A(\cur_mb_mem[198][1] ),
    .B(_06210_),
    .C(_06324_),
    .X(_07029_));
 sky130_fd_sc_hd__and3_1 _11985_ (.A(\cur_mb_mem[82][1] ),
    .B(_06341_),
    .C(_06378_),
    .X(_07030_));
 sky130_fd_sc_hd__and3_1 _11986_ (.A(\cur_mb_mem[152][1] ),
    .B(_06478_),
    .C(_06401_),
    .X(_07031_));
 sky130_fd_sc_hd__a2111o_1 _11987_ (.A1(\cur_mb_mem[65][1] ),
    .A2(_06483_),
    .B1(_07029_),
    .C1(_07030_),
    .D1(_07031_),
    .X(_07032_));
 sky130_fd_sc_hd__and3_1 _11988_ (.A(\cur_mb_mem[165][1] ),
    .B(_06758_),
    .C(_06220_),
    .X(_07033_));
 sky130_fd_sc_hd__and3_1 _11989_ (.A(\cur_mb_mem[67][1] ),
    .B(_06289_),
    .C(_06121_),
    .X(_07034_));
 sky130_fd_sc_hd__and3_1 _11990_ (.A(\cur_mb_mem[178][1] ),
    .B(_06254_),
    .C(_06760_),
    .X(_07035_));
 sky130_fd_sc_hd__a2111o_1 _11991_ (.A1(\cur_mb_mem[74][1] ),
    .A2(_06417_),
    .B1(_07033_),
    .C1(_07034_),
    .D1(_07035_),
    .X(_07036_));
 sky130_fd_sc_hd__and3_1 _11992_ (.A(\cur_mb_mem[106][1] ),
    .B(_05931_),
    .C(_06313_),
    .X(_07037_));
 sky130_fd_sc_hd__and3_1 _11993_ (.A(\cur_mb_mem[121][1] ),
    .B(_06723_),
    .C(_06138_),
    .X(_07038_));
 sky130_fd_sc_hd__and3_1 _11994_ (.A(\cur_mb_mem[123][1] ),
    .B(_06400_),
    .C(_06207_),
    .X(_07039_));
 sky130_fd_sc_hd__a2111o_1 _11995_ (.A1(\cur_mb_mem[41][1] ),
    .A2(_06031_),
    .B1(_07037_),
    .C1(_07038_),
    .D1(_07039_),
    .X(_07040_));
 sky130_fd_sc_hd__and3_1 _11996_ (.A(\cur_mb_mem[169][1] ),
    .B(_06723_),
    .C(_06825_),
    .X(_07041_));
 sky130_fd_sc_hd__and3_2 _11997_ (.A(\cur_mb_mem[20][1] ),
    .B(_06232_),
    .C(_06235_),
    .X(_07042_));
 sky130_fd_sc_hd__and3_2 _11998_ (.A(\cur_mb_mem[213][1] ),
    .B(_06150_),
    .C(_06153_),
    .X(_07043_));
 sky130_fd_sc_hd__a2111o_1 _11999_ (.A1(\cur_mb_mem[112][1] ),
    .A2(_06439_),
    .B1(_07041_),
    .C1(_07042_),
    .D1(_07043_),
    .X(_07044_));
 sky130_fd_sc_hd__or4_2 _12000_ (.A(_07032_),
    .B(_07036_),
    .C(_07040_),
    .D(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__and3_1 _12001_ (.A(\cur_mb_mem[57][1] ),
    .B(_06170_),
    .C(_06038_),
    .X(_07046_));
 sky130_fd_sc_hd__and3_1 _12002_ (.A(\cur_mb_mem[52][1] ),
    .B(_06350_),
    .C(_06744_),
    .X(_07047_));
 sky130_fd_sc_hd__and3_1 _12003_ (.A(\cur_mb_mem[81][1] ),
    .B(_06230_),
    .C(_06841_),
    .X(_07048_));
 sky130_fd_sc_hd__a2111o_1 _12004_ (.A1(\cur_mb_mem[4][1] ),
    .A2(_06162_),
    .B1(_07046_),
    .C1(_07047_),
    .D1(_07048_),
    .X(_07049_));
 sky130_fd_sc_hd__and3_1 _12005_ (.A(\cur_mb_mem[78][1] ),
    .B(_06143_),
    .C(_06046_),
    .X(_07050_));
 sky130_fd_sc_hd__and3_1 _12006_ (.A(\cur_mb_mem[77][1] ),
    .B(_06490_),
    .C(_06121_),
    .X(_07051_));
 sky130_fd_sc_hd__and3_1 _12007_ (.A(\cur_mb_mem[50][1] ),
    .B(_06240_),
    .C(_06254_),
    .X(_07052_));
 sky130_fd_sc_hd__a2111o_1 _12008_ (.A1(\cur_mb_mem[129][1] ),
    .A2(_05966_),
    .B1(_07050_),
    .C1(_07051_),
    .D1(_07052_),
    .X(_07053_));
 sky130_fd_sc_hd__and3_1 _12009_ (.A(\cur_mb_mem[94][1] ),
    .B(_06378_),
    .C(_06435_),
    .X(_07054_));
 sky130_fd_sc_hd__and3_2 _12010_ (.A(\cur_mb_mem[56][1] ),
    .B(_06856_),
    .C(_06455_),
    .X(_07055_));
 sky130_fd_sc_hd__and3_1 _12011_ (.A(\cur_mb_mem[109][1] ),
    .B(_06268_),
    .C(_06762_),
    .X(_07056_));
 sky130_fd_sc_hd__a2111o_2 _12012_ (.A1(\cur_mb_mem[211][1] ),
    .A2(_06349_),
    .B1(_07054_),
    .C1(_07055_),
    .D1(_07056_),
    .X(_07057_));
 sky130_fd_sc_hd__and3_1 _12013_ (.A(\cur_mb_mem[84][1] ),
    .B(_06232_),
    .C(_05914_),
    .X(_07058_));
 sky130_fd_sc_hd__and3_1 _12014_ (.A(\cur_mb_mem[69][1] ),
    .B(_06809_),
    .C(_06208_),
    .X(_07059_));
 sky130_fd_sc_hd__and3_1 _12015_ (.A(\cur_mb_mem[83][1] ),
    .B(_06895_),
    .C(_06980_),
    .X(_07060_));
 sky130_fd_sc_hd__a2111o_1 _12016_ (.A1(\cur_mb_mem[244][1] ),
    .A2(_06167_),
    .B1(_07058_),
    .C1(_07059_),
    .D1(_07060_),
    .X(_07061_));
 sky130_fd_sc_hd__or4_2 _12017_ (.A(_07049_),
    .B(_07053_),
    .C(_07057_),
    .D(_07061_),
    .X(_07062_));
 sky130_fd_sc_hd__and3_2 _12018_ (.A(\cur_mb_mem[219][1] ),
    .B(_06312_),
    .C(_06348_),
    .X(_07063_));
 sky130_fd_sc_hd__and3_1 _12019_ (.A(\cur_mb_mem[73][1] ),
    .B(_06327_),
    .C(_06233_),
    .X(_07064_));
 sky130_fd_sc_hd__and3_2 _12020_ (.A(\cur_mb_mem[205][1] ),
    .B(_06762_),
    .C(_06082_),
    .X(_07065_));
 sky130_fd_sc_hd__a2111o_1 _12021_ (.A1(\cur_mb_mem[1][1] ),
    .A2(_05990_),
    .B1(_07063_),
    .C1(_07064_),
    .D1(_07065_),
    .X(_07066_));
 sky130_fd_sc_hd__and3_1 _12022_ (.A(\cur_mb_mem[164][1] ),
    .B(_06744_),
    .C(_06758_),
    .X(_07067_));
 sky130_fd_sc_hd__and3_1 _12023_ (.A(\cur_mb_mem[214][1] ),
    .B(_06204_),
    .C(_06270_),
    .X(_07068_));
 sky130_fd_sc_hd__and3_1 _12024_ (.A(\cur_mb_mem[171][1] ),
    .B(_06387_),
    .C(_06755_),
    .X(_07069_));
 sky130_fd_sc_hd__a2111o_4 _12025_ (.A1(\cur_mb_mem[209][1] ),
    .A2(_06271_),
    .B1(_07067_),
    .C1(_07068_),
    .D1(_07069_),
    .X(_07070_));
 sky130_fd_sc_hd__and3_1 _12026_ (.A(\cur_mb_mem[5][1] ),
    .B(_06300_),
    .C(_06812_),
    .X(_07071_));
 sky130_fd_sc_hd__and3_1 _12027_ (.A(\cur_mb_mem[97][1] ),
    .B(_05984_),
    .C(_06841_),
    .X(_07072_));
 sky130_fd_sc_hd__and3_4 _12028_ (.A(\cur_mb_mem[203][1] ),
    .B(_06387_),
    .C(_06967_),
    .X(_07073_));
 sky130_fd_sc_hd__a2111o_1 _12029_ (.A1(\cur_mb_mem[66][1] ),
    .A2(_06368_),
    .B1(_07071_),
    .C1(_07072_),
    .D1(_07073_),
    .X(_07074_));
 sky130_fd_sc_hd__buf_12 _12030_ (.A(_05952_),
    .X(_07075_));
 sky130_fd_sc_hd__and3_1 _12031_ (.A(\cur_mb_mem[222][1] ),
    .B(_06814_),
    .C(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__and3_1 _12032_ (.A(\cur_mb_mem[173][1] ),
    .B(_06056_),
    .C(_06192_),
    .X(_07077_));
 sky130_fd_sc_hd__buf_6 _12033_ (.A(_06050_),
    .X(_07078_));
 sky130_fd_sc_hd__and3_1 _12034_ (.A(\cur_mb_mem[125][1] ),
    .B(_06246_),
    .C(_07078_),
    .X(_07079_));
 sky130_fd_sc_hd__a2111o_2 _12035_ (.A1(\cur_mb_mem[19][1] ),
    .A2(_06282_),
    .B1(_07076_),
    .C1(_07077_),
    .D1(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__or4_2 _12036_ (.A(_07066_),
    .B(_07070_),
    .C(_07074_),
    .D(_07080_),
    .X(_07081_));
 sky130_fd_sc_hd__and3_1 _12037_ (.A(\cur_mb_mem[13][1] ),
    .B(_06202_),
    .C(_06490_),
    .X(_07082_));
 sky130_fd_sc_hd__and3_2 _12038_ (.A(\cur_mb_mem[240][1] ),
    .B(_06916_),
    .C(_06772_),
    .X(_07083_));
 sky130_fd_sc_hd__clkbuf_16 _12039_ (.A(_05953_),
    .X(_07084_));
 sky130_fd_sc_hd__and3_1 _12040_ (.A(\cur_mb_mem[174][1] ),
    .B(_07084_),
    .C(_07001_),
    .X(_07085_));
 sky130_fd_sc_hd__a2111o_1 _12041_ (.A1(\cur_mb_mem[22][1] ),
    .A2(_06242_),
    .B1(_07082_),
    .C1(_07083_),
    .D1(_07085_),
    .X(_07086_));
 sky130_fd_sc_hd__and3_2 _12042_ (.A(\cur_mb_mem[202][1] ),
    .B(_06442_),
    .C(_06789_),
    .X(_07087_));
 sky130_fd_sc_hd__and3_1 _12043_ (.A(\cur_mb_mem[241][1] ),
    .B(_06032_),
    .C(net227),
    .X(_07088_));
 sky130_fd_sc_hd__and3_2 _12044_ (.A(\cur_mb_mem[75][1] ),
    .B(_05917_),
    .C(_06022_),
    .X(_07089_));
 sky130_fd_sc_hd__and3_1 _12045_ (.A(\cur_mb_mem[186][1] ),
    .B(_05931_),
    .C(_06013_),
    .X(_07090_));
 sky130_fd_sc_hd__or4_1 _12046_ (.A(_07087_),
    .B(_07088_),
    .C(_07089_),
    .D(_07090_),
    .X(_07091_));
 sky130_fd_sc_hd__and3_1 _12047_ (.A(\cur_mb_mem[245][1] ),
    .B(_06165_),
    .C(_06208_),
    .X(_07092_));
 sky130_fd_sc_hd__and3_1 _12048_ (.A(\cur_mb_mem[196][1] ),
    .B(_06215_),
    .C(_06967_),
    .X(_07093_));
 sky130_fd_sc_hd__and3_1 _12049_ (.A(\cur_mb_mem[160][1] ),
    .B(_07001_),
    .C(_06315_),
    .X(_07094_));
 sky130_fd_sc_hd__a2111o_1 _12050_ (.A1(\cur_mb_mem[101][1] ),
    .A2(_06269_),
    .B1(_07092_),
    .C1(_07093_),
    .D1(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__buf_12 _12051_ (.A(net252),
    .X(_07096_));
 sky130_fd_sc_hd__and3_1 _12052_ (.A(\cur_mb_mem[6][1] ),
    .B(_07096_),
    .C(_06191_),
    .X(_07097_));
 sky130_fd_sc_hd__and3_1 _12053_ (.A(\cur_mb_mem[208][1] ),
    .B(_05947_),
    .C(_06748_),
    .X(_07098_));
 sky130_fd_sc_hd__buf_6 _12054_ (.A(_06079_),
    .X(_07099_));
 sky130_fd_sc_hd__buf_4 _12055_ (.A(_05977_),
    .X(_07100_));
 sky130_fd_sc_hd__and3_1 _12056_ (.A(\cur_mb_mem[146][1] ),
    .B(_07099_),
    .C(_07100_),
    .X(_07101_));
 sky130_fd_sc_hd__a2111o_2 _12057_ (.A1(\cur_mb_mem[166][1] ),
    .A2(_06193_),
    .B1(_07097_),
    .C1(_07098_),
    .D1(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__or4_2 _12058_ (.A(_07086_),
    .B(_07091_),
    .C(_07095_),
    .D(_07102_),
    .X(_07103_));
 sky130_fd_sc_hd__or4_1 _12059_ (.A(_07045_),
    .B(_07062_),
    .C(_07081_),
    .D(_07103_),
    .X(_07104_));
 sky130_fd_sc_hd__a32o_1 _12060_ (.A1(\cur_mb_mem[224][1] ),
    .A2(_05971_),
    .A3(_06224_),
    .B1(_06305_),
    .B2(\cur_mb_mem[143][1] ),
    .X(_07105_));
 sky130_fd_sc_hd__a32o_1 _12061_ (.A1(\cur_mb_mem[230][1] ),
    .A2(_06186_),
    .A3(_06224_),
    .B1(_06069_),
    .B2(\cur_mb_mem[111][1] ),
    .X(_07106_));
 sky130_fd_sc_hd__a2111o_1 _12062_ (.A1(\cur_mb_mem[127][1] ),
    .A2(_06101_),
    .B1(_07105_),
    .C1(_07106_),
    .D1(_06185_),
    .X(_07107_));
 sky130_fd_sc_hd__and3_1 _12063_ (.A(\cur_mb_mem[18][1] ),
    .B(_06079_),
    .C(_05974_),
    .X(_07108_));
 sky130_fd_sc_hd__and3_1 _12064_ (.A(\cur_mb_mem[44][1] ),
    .B(_05901_),
    .C(_06005_),
    .X(_07109_));
 sky130_fd_sc_hd__and3_2 _12065_ (.A(\cur_mb_mem[227][1] ),
    .B(_06061_),
    .C(_05997_),
    .X(_07110_));
 sky130_fd_sc_hd__and3_1 _12066_ (.A(\cur_mb_mem[36][1] ),
    .B(_06026_),
    .C(_06005_),
    .X(_07111_));
 sky130_fd_sc_hd__or4_2 _12067_ (.A(_07108_),
    .B(_07109_),
    .C(_07110_),
    .D(_07111_),
    .X(_07112_));
 sky130_fd_sc_hd__and3_1 _12068_ (.A(\cur_mb_mem[228][1] ),
    .B(_06026_),
    .C(_06116_),
    .X(_07113_));
 sky130_fd_sc_hd__and3_2 _12069_ (.A(\cur_mb_mem[79][1] ),
    .B(_06120_),
    .C(_06233_),
    .X(_07114_));
 sky130_fd_sc_hd__and3_1 _12070_ (.A(\cur_mb_mem[234][1] ),
    .B(_05957_),
    .C(_06766_),
    .X(_07115_));
 sky130_fd_sc_hd__a2111o_1 _12071_ (.A1(\cur_mb_mem[15][1] ),
    .A2(_06295_),
    .B1(_07113_),
    .C1(_07114_),
    .D1(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__and3_1 _12072_ (.A(\cur_mb_mem[49][1] ),
    .B(_06350_),
    .C(_05995_),
    .X(_07117_));
 sky130_fd_sc_hd__and3_1 _12073_ (.A(\cur_mb_mem[48][1] ),
    .B(_06856_),
    .C(_06815_),
    .X(_07118_));
 sky130_fd_sc_hd__and3_1 _12074_ (.A(\cur_mb_mem[62][1] ),
    .B(_06198_),
    .C(_07075_),
    .X(_07119_));
 sky130_fd_sc_hd__a2111o_4 _12075_ (.A1(\cur_mb_mem[25][1] ),
    .A2(_06489_),
    .B1(_07117_),
    .C1(_07118_),
    .D1(_07119_),
    .X(_07120_));
 sky130_fd_sc_hd__and3_1 _12076_ (.A(\cur_mb_mem[63][1] ),
    .B(_06466_),
    .C(_06856_),
    .X(_07121_));
 sky130_fd_sc_hd__and3_1 _12077_ (.A(\cur_mb_mem[239][1] ),
    .B(_06149_),
    .C(_06247_),
    .X(_07122_));
 sky130_fd_sc_hd__and3_1 _12078_ (.A(\cur_mb_mem[90][1] ),
    .B(_05905_),
    .C(_06895_),
    .X(_07123_));
 sky130_fd_sc_hd__a2111o_1 _12079_ (.A1(\cur_mb_mem[191][1] ),
    .A2(_06467_),
    .B1(_07121_),
    .C1(_07122_),
    .D1(_07123_),
    .X(_07124_));
 sky130_fd_sc_hd__or4_2 _12080_ (.A(_07112_),
    .B(_07116_),
    .C(_07120_),
    .D(_07124_),
    .X(_07125_));
 sky130_fd_sc_hd__a32o_1 _12081_ (.A1(\cur_mb_mem[218][1] ),
    .A2(_05958_),
    .A3(_05948_),
    .B1(_06487_),
    .B2(\cur_mb_mem[142][1] ),
    .X(_07126_));
 sky130_fd_sc_hd__a32o_1 _12082_ (.A1(\cur_mb_mem[105][1] ),
    .A2(_05910_),
    .A3(_06298_),
    .B1(_06034_),
    .B2(\cur_mb_mem[253][1] ),
    .X(_07127_));
 sky130_fd_sc_hd__or2_2 _12083_ (.A(_07126_),
    .B(_07127_),
    .X(_07128_));
 sky130_fd_sc_hd__a32o_1 _12084_ (.A1(\cur_mb_mem[251][1] ),
    .A2(_04430_),
    .A3(_06261_),
    .B1(_06414_),
    .B2(\cur_mb_mem[102][1] ),
    .X(_07129_));
 sky130_fd_sc_hd__a22o_2 _12085_ (.A1(\cur_mb_mem[180][1] ),
    .A2(_06217_),
    .B1(_06234_),
    .B2(\cur_mb_mem[68][1] ),
    .X(_07130_));
 sky130_fd_sc_hd__and3_1 _12086_ (.A(\cur_mb_mem[117][1] ),
    .B(_06207_),
    .C(_06208_),
    .X(_07131_));
 sky130_fd_sc_hd__and3_1 _12087_ (.A(\cur_mb_mem[201][1] ),
    .B(_06903_),
    .C(_06967_),
    .X(_07132_));
 sky130_fd_sc_hd__and3_2 _12088_ (.A(\cur_mb_mem[136][1] ),
    .B(_06774_),
    .C(_06859_),
    .X(_07133_));
 sky130_fd_sc_hd__a2111o_1 _12089_ (.A1(\cur_mb_mem[158][1] ),
    .A2(_06436_),
    .B1(_07131_),
    .C1(_07132_),
    .D1(_07133_),
    .X(_07134_));
 sky130_fd_sc_hd__and3_1 _12090_ (.A(\cur_mb_mem[212][1] ),
    .B(_06215_),
    .C(_06150_),
    .X(_07135_));
 sky130_fd_sc_hd__and3_1 _12091_ (.A(\cur_mb_mem[192][1] ),
    .B(_06997_),
    .C(_06315_),
    .X(_07136_));
 sky130_fd_sc_hd__buf_6 _12092_ (.A(_04429_),
    .X(_07137_));
 sky130_fd_sc_hd__and3_1 _12093_ (.A(\cur_mb_mem[252][1] ),
    .B(_07137_),
    .C(_06920_),
    .X(_07138_));
 sky130_fd_sc_hd__a2111o_1 _12094_ (.A1(\cur_mb_mem[145][1] ),
    .A2(_06252_),
    .B1(_07135_),
    .C1(_07136_),
    .D1(_07138_),
    .X(_07139_));
 sky130_fd_sc_hd__or4_2 _12095_ (.A(_07129_),
    .B(_07130_),
    .C(_07134_),
    .D(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__or4_2 _12096_ (.A(_07107_),
    .B(_07125_),
    .C(_07128_),
    .D(_07140_),
    .X(_07141_));
 sky130_fd_sc_hd__and3_1 _12097_ (.A(\cur_mb_mem[148][1] ),
    .B(_06744_),
    .C(_06434_),
    .X(_07142_));
 sky130_fd_sc_hd__and3_1 _12098_ (.A(\cur_mb_mem[92][1] ),
    .B(_06718_),
    .C(_06931_),
    .X(_07143_));
 sky130_fd_sc_hd__and3_1 _12099_ (.A(\cur_mb_mem[122][1] ),
    .B(_06960_),
    .C(_06207_),
    .X(_07144_));
 sky130_fd_sc_hd__a2111o_1 _12100_ (.A1(\cur_mb_mem[179][1] ),
    .A2(_06356_),
    .B1(_07142_),
    .C1(_07143_),
    .D1(_07144_),
    .X(_07145_));
 sky130_fd_sc_hd__and3_1 _12101_ (.A(\cur_mb_mem[140][1] ),
    .B(_06718_),
    .C(_06382_),
    .X(_07146_));
 sky130_fd_sc_hd__and3_2 _12102_ (.A(\cur_mb_mem[54][1] ),
    .B(_06856_),
    .C(_06204_),
    .X(_07147_));
 sky130_fd_sc_hd__and3_1 _12103_ (.A(\cur_mb_mem[181][1] ),
    .B(_06830_),
    .C(_06208_),
    .X(_07148_));
 sky130_fd_sc_hd__a2111o_1 _12104_ (.A1(\cur_mb_mem[14][1] ),
    .A2(_06367_),
    .B1(_07146_),
    .C1(_07147_),
    .D1(_07148_),
    .X(_07149_));
 sky130_fd_sc_hd__and3_1 _12105_ (.A(\cur_mb_mem[221][1] ),
    .B(_06490_),
    .C(_06270_),
    .X(_07150_));
 sky130_fd_sc_hd__and3_1 _12106_ (.A(\cur_mb_mem[124][1] ),
    .B(_06754_),
    .C(_06138_),
    .X(_07151_));
 sky130_fd_sc_hd__and3_1 _12107_ (.A(\cur_mb_mem[9][1] ),
    .B(_07096_),
    .C(_06903_),
    .X(_07152_));
 sky130_fd_sc_hd__a2111o_2 _12108_ (.A1(\cur_mb_mem[27][1] ),
    .A2(_06476_),
    .B1(_07150_),
    .C1(_07151_),
    .D1(_07152_),
    .X(_07153_));
 sky130_fd_sc_hd__and3_1 _12109_ (.A(\cur_mb_mem[16][1] ),
    .B(_05970_),
    .C(_06235_),
    .X(_07154_));
 sky130_fd_sc_hd__and3_1 _12110_ (.A(\cur_mb_mem[188][1] ),
    .B(_06937_),
    .C(_06830_),
    .X(_07155_));
 sky130_fd_sc_hd__and3_1 _12111_ (.A(\cur_mb_mem[72][1] ),
    .B(_06832_),
    .C(_06023_),
    .X(_07156_));
 sky130_fd_sc_hd__a2111o_1 _12112_ (.A1(\cur_mb_mem[40][1] ),
    .A2(_06485_),
    .B1(_07154_),
    .C1(_07155_),
    .D1(_07156_),
    .X(_07157_));
 sky130_fd_sc_hd__or4_1 _12113_ (.A(_07145_),
    .B(_07149_),
    .C(_07153_),
    .D(_07157_),
    .X(_07158_));
 sky130_fd_sc_hd__and3_2 _12114_ (.A(\cur_mb_mem[131][1] ),
    .B(_06355_),
    .C(_06382_),
    .X(_07159_));
 sky130_fd_sc_hd__and3_1 _12115_ (.A(\cur_mb_mem[130][1] ),
    .B(_06254_),
    .C(_06842_),
    .X(_07160_));
 sky130_fd_sc_hd__and3_2 _12116_ (.A(\cur_mb_mem[120][1] ),
    .B(_05982_),
    .C(_06207_),
    .X(_07161_));
 sky130_fd_sc_hd__a2111o_1 _12117_ (.A1(\cur_mb_mem[12][1] ),
    .A2(_05928_),
    .B1(_07159_),
    .C1(_07160_),
    .D1(_07161_),
    .X(_07162_));
 sky130_fd_sc_hd__and3_1 _12118_ (.A(\cur_mb_mem[217][1] ),
    .B(_06327_),
    .C(_06270_),
    .X(_07163_));
 sky130_fd_sc_hd__and3_1 _12119_ (.A(\cur_mb_mem[155][1] ),
    .B(_06474_),
    .C(_06401_),
    .X(_07164_));
 sky130_fd_sc_hd__and3_1 _12120_ (.A(\cur_mb_mem[149][1] ),
    .B(_06747_),
    .C(_06794_),
    .X(_07165_));
 sky130_fd_sc_hd__a2111o_2 _12121_ (.A1(\cur_mb_mem[11][1] ),
    .A2(_06301_),
    .B1(_07163_),
    .C1(_07164_),
    .D1(_07165_),
    .X(_07166_));
 sky130_fd_sc_hd__and3_1 _12122_ (.A(\cur_mb_mem[100][1] ),
    .B(_06166_),
    .C(_06045_),
    .X(_07167_));
 sky130_fd_sc_hd__and3_1 _12123_ (.A(\cur_mb_mem[133][1] ),
    .B(_06842_),
    .C(_06147_),
    .X(_07168_));
 sky130_fd_sc_hd__and3_1 _12124_ (.A(\cur_mb_mem[76][1] ),
    .B(_06937_),
    .C(_06057_),
    .X(_07169_));
 sky130_fd_sc_hd__a2111o_1 _12125_ (.A1(\cur_mb_mem[184][1] ),
    .A2(_06479_),
    .B1(_07167_),
    .C1(_07168_),
    .D1(_07169_),
    .X(_07170_));
 sky130_fd_sc_hd__and3_1 _12126_ (.A(\cur_mb_mem[176][1] ),
    .B(_06830_),
    .C(_06772_),
    .X(_07171_));
 sky130_fd_sc_hd__and3_1 _12127_ (.A(\cur_mb_mem[88][1] ),
    .B(_06832_),
    .C(_06927_),
    .X(_07172_));
 sky130_fd_sc_hd__and3_1 _12128_ (.A(\cur_mb_mem[86][1] ),
    .B(_06895_),
    .C(_06191_),
    .X(_07173_));
 sky130_fd_sc_hd__a2111o_1 _12129_ (.A1(\cur_mb_mem[182][1] ),
    .A2(_06205_),
    .B1(_07171_),
    .C1(_07172_),
    .D1(_07173_),
    .X(_07174_));
 sky130_fd_sc_hd__or4_1 _12130_ (.A(_07162_),
    .B(_07166_),
    .C(_07170_),
    .D(_07174_),
    .X(_07175_));
 sky130_fd_sc_hd__and3_1 _12131_ (.A(\cur_mb_mem[108][1] ),
    .B(_06718_),
    .C(_06045_),
    .X(_07176_));
 sky130_fd_sc_hd__and3_1 _12132_ (.A(\cur_mb_mem[132][1] ),
    .B(_06232_),
    .C(_06842_),
    .X(_07177_));
 sky130_fd_sc_hd__and3_1 _12133_ (.A(\cur_mb_mem[163][1] ),
    .B(_06980_),
    .C(_06192_),
    .X(_07178_));
 sky130_fd_sc_hd__a2111o_1 _12134_ (.A1(\cur_mb_mem[3][1] ),
    .A2(_06290_),
    .B1(_07176_),
    .C1(_07177_),
    .D1(_07178_),
    .X(_07179_));
 sky130_fd_sc_hd__and3_1 _12135_ (.A(\cur_mb_mem[197][1] ),
    .B(_06352_),
    .C(_06812_),
    .X(_07180_));
 sky130_fd_sc_hd__and3_1 _12136_ (.A(\cur_mb_mem[195][1] ),
    .B(_06770_),
    .C(_06352_),
    .X(_07181_));
 sky130_fd_sc_hd__and3_2 _12137_ (.A(\cur_mb_mem[89][1] ),
    .B(_06834_),
    .C(_06927_),
    .X(_07182_));
 sky130_fd_sc_hd__a2111o_2 _12138_ (.A1(\cur_mb_mem[10][1] ),
    .A2(_06408_),
    .B1(_07180_),
    .C1(_07181_),
    .D1(_07182_),
    .X(_07183_));
 sky130_fd_sc_hd__and3_1 _12139_ (.A(\cur_mb_mem[144][1] ),
    .B(_06401_),
    .C(_05970_),
    .X(_07184_));
 sky130_fd_sc_hd__and3_2 _12140_ (.A(\cur_mb_mem[206][1] ),
    .B(_07075_),
    .C(_06082_),
    .X(_07185_));
 sky130_fd_sc_hd__and3_1 _12141_ (.A(\cur_mb_mem[150][1] ),
    .B(_06191_),
    .C(_06152_),
    .X(_07186_));
 sky130_fd_sc_hd__a2111o_1 _12142_ (.A1(\cur_mb_mem[21][1] ),
    .A2(_06236_),
    .B1(_07184_),
    .C1(_07185_),
    .D1(_07186_),
    .X(_07187_));
 sky130_fd_sc_hd__and3_1 _12143_ (.A(\cur_mb_mem[32][1] ),
    .B(_06952_),
    .C(_06772_),
    .X(_07188_));
 sky130_fd_sc_hd__and3_1 _12144_ (.A(\cur_mb_mem[137][1] ),
    .B(_06834_),
    .C(_06859_),
    .X(_07189_));
 sky130_fd_sc_hd__and3_1 _12145_ (.A(\cur_mb_mem[33][1] ),
    .B(_06044_),
    .C(_05993_),
    .X(_07190_));
 sky130_fd_sc_hd__a2111o_1 _12146_ (.A1(\cur_mb_mem[193][1] ),
    .A2(_06354_),
    .B1(_07188_),
    .C1(_07189_),
    .D1(_07190_),
    .X(_07191_));
 sky130_fd_sc_hd__or4_1 _12147_ (.A(_07179_),
    .B(_07183_),
    .C(_07187_),
    .D(_07191_),
    .X(_07192_));
 sky130_fd_sc_hd__and3_1 _12148_ (.A(\cur_mb_mem[38][1] ),
    .B(_06343_),
    .C(_06199_),
    .X(_07193_));
 sky130_fd_sc_hd__and3_2 _12149_ (.A(\cur_mb_mem[147][1] ),
    .B(_06770_),
    .C(_06747_),
    .X(_07194_));
 sky130_fd_sc_hd__buf_4 _12150_ (.A(_06851_),
    .X(_07195_));
 sky130_fd_sc_hd__and3_1 _12151_ (.A(\cur_mb_mem[119][1] ),
    .B(_07078_),
    .C(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__a2111o_1 _12152_ (.A1(\cur_mb_mem[210][1] ),
    .A2(_06342_),
    .B1(_07193_),
    .C1(_07194_),
    .D1(_07196_),
    .X(_07197_));
 sky130_fd_sc_hd__and3_1 _12153_ (.A(\cur_mb_mem[135][1] ),
    .B(_06708_),
    .C(_06842_),
    .X(_07198_));
 sky130_fd_sc_hd__and3_1 _12154_ (.A(\cur_mb_mem[103][1] ),
    .B(_06268_),
    .C(_06896_),
    .X(_07199_));
 sky130_fd_sc_hd__and3_1 _12155_ (.A(\cur_mb_mem[183][1] ),
    .B(_06877_),
    .C(_07195_),
    .X(_07200_));
 sky130_fd_sc_hd__a2111o_1 _12156_ (.A1(\cur_mb_mem[71][1] ),
    .A2(_06460_),
    .B1(_07198_),
    .C1(_07199_),
    .D1(_07200_),
    .X(_07201_));
 sky130_fd_sc_hd__and3_2 _12157_ (.A(\cur_mb_mem[141][1] ),
    .B(_06056_),
    .C(_06146_),
    .X(_07202_));
 sky130_fd_sc_hd__and3_1 _12158_ (.A(\cur_mb_mem[46][1] ),
    .B(_06087_),
    .C(_06000_),
    .X(_07203_));
 sky130_fd_sc_hd__and3_1 _12159_ (.A(\cur_mb_mem[177][1] ),
    .B(_06216_),
    .C(_05993_),
    .X(_07204_));
 sky130_fd_sc_hd__a2111o_1 _12160_ (.A1(\cur_mb_mem[134][1] ),
    .A2(_06211_),
    .B1(_07202_),
    .C1(_07203_),
    .D1(_07204_),
    .X(_07205_));
 sky130_fd_sc_hd__and3_1 _12161_ (.A(\cur_mb_mem[23][1] ),
    .B(_07195_),
    .C(_06001_),
    .X(_07206_));
 sky130_fd_sc_hd__and3_2 _12162_ (.A(\cur_mb_mem[207][1] ),
    .B(_04423_),
    .C(_06997_),
    .X(_07207_));
 sky130_fd_sc_hd__and3_1 _12163_ (.A(\cur_mb_mem[128][1] ),
    .B(_06315_),
    .C(_05935_),
    .X(_07208_));
 sky130_fd_sc_hd__a2111o_1 _12164_ (.A1(\cur_mb_mem[61][1] ),
    .A2(_06359_),
    .B1(_07206_),
    .C1(_07207_),
    .D1(_07208_),
    .X(_07209_));
 sky130_fd_sc_hd__or4_2 _12165_ (.A(_07197_),
    .B(_07201_),
    .C(_07205_),
    .D(_07209_),
    .X(_07210_));
 sky130_fd_sc_hd__or4_2 _12166_ (.A(_07158_),
    .B(_07175_),
    .C(_07192_),
    .D(_07210_),
    .X(_07211_));
 sky130_fd_sc_hd__and3_1 _12167_ (.A(\cur_mb_mem[236][1] ),
    .B(_06754_),
    .C(_06255_),
    .X(_07212_));
 sky130_fd_sc_hd__and3_1 _12168_ (.A(\cur_mb_mem[255][1] ),
    .B(_06466_),
    .C(_06916_),
    .X(_07213_));
 sky130_fd_sc_hd__and3_2 _12169_ (.A(\cur_mb_mem[151][1] ),
    .B(_06152_),
    .C(_06896_),
    .X(_07214_));
 sky130_fd_sc_hd__a2111o_1 _12170_ (.A1(\cur_mb_mem[231][1] ),
    .A2(_06180_),
    .B1(_07212_),
    .C1(_07213_),
    .D1(_07214_),
    .X(_07215_));
 sky130_fd_sc_hd__and3_1 _12171_ (.A(\cur_mb_mem[7][1] ),
    .B(_06202_),
    .C(_06372_),
    .X(_07216_));
 sky130_fd_sc_hd__and3_1 _12172_ (.A(\cur_mb_mem[235][1] ),
    .B(_06400_),
    .C(_06247_),
    .X(_07217_));
 sky130_fd_sc_hd__and3_1 _12173_ (.A(\cur_mb_mem[167][1] ),
    .B(_07001_),
    .C(_06896_),
    .X(_07218_));
 sky130_fd_sc_hd__a2111o_1 _12174_ (.A1(\cur_mb_mem[226][1] ),
    .A2(_06256_),
    .B1(_07216_),
    .C1(_07217_),
    .D1(_07218_),
    .X(_07219_));
 sky130_fd_sc_hd__and3_1 _12175_ (.A(\cur_mb_mem[91][1] ),
    .B(_06400_),
    .C(_06230_),
    .X(_07220_));
 sky130_fd_sc_hd__and3_1 _12176_ (.A(\cur_mb_mem[45][1] ),
    .B(_06952_),
    .C(_06056_),
    .X(_07221_));
 sky130_fd_sc_hd__and3_1 _12177_ (.A(\cur_mb_mem[242][1] ),
    .B(_07137_),
    .C(_06380_),
    .X(_07222_));
 sky130_fd_sc_hd__a2111o_4 _12178_ (.A1(\cur_mb_mem[194][1] ),
    .A2(_06083_),
    .B1(_07220_),
    .C1(_07221_),
    .D1(_07222_),
    .X(_07223_));
 sky130_fd_sc_hd__and3_1 _12179_ (.A(\cur_mb_mem[233][1] ),
    .B(_06834_),
    .C(_06247_),
    .X(_07224_));
 sky130_fd_sc_hd__and3_1 _12180_ (.A(\cur_mb_mem[232][1] ),
    .B(_06832_),
    .C(_06775_),
    .X(_07225_));
 sky130_fd_sc_hd__and3_1 _12181_ (.A(\cur_mb_mem[189][1] ),
    .B(_06246_),
    .C(_06216_),
    .X(_07226_));
 sky130_fd_sc_hd__a2111o_1 _12182_ (.A1(\cur_mb_mem[35][1] ),
    .A2(_06088_),
    .B1(_07224_),
    .C1(_07225_),
    .D1(_07226_),
    .X(_07227_));
 sky130_fd_sc_hd__or4_2 _12183_ (.A(_07215_),
    .B(_07219_),
    .C(_07223_),
    .D(_07227_),
    .X(_07228_));
 sky130_fd_sc_hd__and3_1 _12184_ (.A(\cur_mb_mem[199][1] ),
    .B(_06352_),
    .C(_06372_),
    .X(_07229_));
 sky130_fd_sc_hd__and3_1 _12185_ (.A(\cur_mb_mem[175][1] ),
    .B(_06149_),
    .C(_06755_),
    .X(_07230_));
 sky130_fd_sc_hd__and3_1 _12186_ (.A(\cur_mb_mem[87][1] ),
    .B(_06895_),
    .C(_06896_),
    .X(_07231_));
 sky130_fd_sc_hd__a2111o_1 _12187_ (.A1(\cur_mb_mem[215][1] ),
    .A2(_06447_),
    .B1(_07229_),
    .C1(_07230_),
    .D1(_07231_),
    .X(_07232_));
 sky130_fd_sc_hd__and3_1 _12188_ (.A(\cur_mb_mem[238][1] ),
    .B(_07075_),
    .C(_06766_),
    .X(_07233_));
 sky130_fd_sc_hd__and3_1 _12189_ (.A(\cur_mb_mem[47][1] ),
    .B(_06149_),
    .C(_06952_),
    .X(_07234_));
 sky130_fd_sc_hd__buf_6 _12190_ (.A(_06849_),
    .X(_07235_));
 sky130_fd_sc_hd__and3_1 _12191_ (.A(\cur_mb_mem[55][1] ),
    .B(_07235_),
    .C(_07195_),
    .X(_07236_));
 sky130_fd_sc_hd__a2111o_1 _12192_ (.A1(\cur_mb_mem[37][1] ),
    .A2(_06344_),
    .B1(_07233_),
    .C1(_07234_),
    .D1(_07236_),
    .X(_07237_));
 sky130_fd_sc_hd__and3_1 _12193_ (.A(\cur_mb_mem[162][1] ),
    .B(_06080_),
    .C(_06755_),
    .X(_07238_));
 sky130_fd_sc_hd__and3_2 _12194_ (.A(\cur_mb_mem[114][1] ),
    .B(_06908_),
    .C(_07078_),
    .X(_07239_));
 sky130_fd_sc_hd__and3_1 _12195_ (.A(\cur_mb_mem[60][1] ),
    .B(_07235_),
    .C(_05902_),
    .X(_07240_));
 sky130_fd_sc_hd__a2111o_1 _12196_ (.A1(\cur_mb_mem[34][1] ),
    .A2(_06393_),
    .B1(_07238_),
    .C1(_07239_),
    .D1(_07240_),
    .X(_07241_));
 sky130_fd_sc_hd__and3_1 _12197_ (.A(\cur_mb_mem[229][1] ),
    .B(_06153_),
    .C(_06918_),
    .X(_07242_));
 sky130_fd_sc_hd__and3_1 _12198_ (.A(\cur_mb_mem[39][1] ),
    .B(_06044_),
    .C(_07195_),
    .X(_07243_));
 sky130_fd_sc_hd__and3_1 _12199_ (.A(\cur_mb_mem[243][1] ),
    .B(_07137_),
    .C(_06086_),
    .X(_07244_));
 sky130_fd_sc_hd__a2111o_2 _12200_ (.A1(\cur_mb_mem[237][1] ),
    .A2(_06248_),
    .B1(_07242_),
    .C1(_07243_),
    .D1(_07244_),
    .X(_07245_));
 sky130_fd_sc_hd__or4_1 _12201_ (.A(_07232_),
    .B(_07237_),
    .C(_07241_),
    .D(_07245_),
    .X(_07246_));
 sky130_fd_sc_hd__and3_1 _12202_ (.A(\cur_mb_mem[107][1] ),
    .B(_06400_),
    .C(_05984_),
    .X(_07247_));
 sky130_fd_sc_hd__and3_1 _12203_ (.A(\cur_mb_mem[138][1] ),
    .B(_06960_),
    .C(_06146_),
    .X(_07248_));
 sky130_fd_sc_hd__and3_1 _12204_ (.A(\cur_mb_mem[156][1] ),
    .B(_05902_),
    .C(_07100_),
    .X(_07249_));
 sky130_fd_sc_hd__a2111o_2 _12205_ (.A1(\cur_mb_mem[70][1] ),
    .A2(_06144_),
    .B1(_07247_),
    .C1(_07248_),
    .D1(_07249_),
    .X(_07250_));
 sky130_fd_sc_hd__and3_4 _12206_ (.A(\cur_mb_mem[225][1] ),
    .B(_06912_),
    .C(_06766_),
    .X(_07251_));
 sky130_fd_sc_hd__and3_1 _12207_ (.A(\cur_mb_mem[247][1] ),
    .B(_06902_),
    .C(_06708_),
    .X(_07252_));
 sky130_fd_sc_hd__buf_8 _12208_ (.A(_06050_),
    .X(_07253_));
 sky130_fd_sc_hd__and3_1 _12209_ (.A(\cur_mb_mem[115][1] ),
    .B(_06086_),
    .C(_07253_),
    .X(_07254_));
 sky130_fd_sc_hd__a2111o_1 _12210_ (.A1(\cur_mb_mem[43][1] ),
    .A2(_06006_),
    .B1(_07251_),
    .C1(_07252_),
    .D1(_07254_),
    .X(_07255_));
 sky130_fd_sc_hd__and3_2 _12211_ (.A(\cur_mb_mem[2][1] ),
    .B(_06707_),
    .C(_06080_),
    .X(_07256_));
 sky130_fd_sc_hd__and3_4 _12212_ (.A(\cur_mb_mem[51][1] ),
    .B(_07235_),
    .C(_06980_),
    .X(_07257_));
 sky130_fd_sc_hd__and3_1 _12213_ (.A(\cur_mb_mem[96][1] ),
    .B(_06413_),
    .C(_06315_),
    .X(_07258_));
 sky130_fd_sc_hd__a2111o_2 _12214_ (.A1(\cur_mb_mem[104][1] ),
    .A2(_05985_),
    .B1(_07256_),
    .C1(_07257_),
    .D1(_07258_),
    .X(_07259_));
 sky130_fd_sc_hd__and3_1 _12215_ (.A(\cur_mb_mem[220][1] ),
    .B(_05902_),
    .C(_05947_),
    .X(_07260_));
 sky130_fd_sc_hd__and3_1 _12216_ (.A(\cur_mb_mem[187][1] ),
    .B(_06942_),
    .C(_06216_),
    .X(_07261_));
 sky130_fd_sc_hd__and3_1 _12217_ (.A(\cur_mb_mem[126][1] ),
    .B(_07021_),
    .C(_05954_),
    .X(_07262_));
 sky130_fd_sc_hd__a2111o_1 _12218_ (.A1(\cur_mb_mem[139][1] ),
    .A2(_06388_),
    .B1(_07260_),
    .C1(_07261_),
    .D1(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__or4_2 _12219_ (.A(_07250_),
    .B(_07255_),
    .C(_07259_),
    .D(_07263_),
    .X(_07264_));
 sky130_fd_sc_hd__and3_1 _12220_ (.A(\cur_mb_mem[17][1] ),
    .B(_06251_),
    .C(_06001_),
    .X(_07265_));
 sky130_fd_sc_hd__and3_2 _12221_ (.A(\cur_mb_mem[64][1] ),
    .B(_06057_),
    .C(_06748_),
    .X(_07266_));
 sky130_fd_sc_hd__and3_1 _12222_ (.A(\cur_mb_mem[118][1] ),
    .B(_07021_),
    .C(_06186_),
    .X(_07267_));
 sky130_fd_sc_hd__a2111o_1 _12223_ (.A1(\cur_mb_mem[85][1] ),
    .A2(_06231_),
    .B1(_07265_),
    .C1(_07266_),
    .D1(_07267_),
    .X(_07268_));
 sky130_fd_sc_hd__and3_1 _12224_ (.A(\cur_mb_mem[58][1] ),
    .B(_07235_),
    .C(_06960_),
    .X(_07269_));
 sky130_fd_sc_hd__and3_1 _12225_ (.A(\cur_mb_mem[59][1] ),
    .B(_07235_),
    .C(_06942_),
    .X(_07270_));
 sky130_fd_sc_hd__and3_2 _12226_ (.A(\cur_mb_mem[157][1] ),
    .B(_05945_),
    .C(_07100_),
    .X(_07271_));
 sky130_fd_sc_hd__a2111o_1 _12227_ (.A1(\cur_mb_mem[161][1] ),
    .A2(_06334_),
    .B1(_07269_),
    .C1(_07270_),
    .D1(_07271_),
    .X(_07272_));
 sky130_fd_sc_hd__and3_1 _12228_ (.A(\cur_mb_mem[204][1] ),
    .B(_05902_),
    .C(_06997_),
    .X(_07273_));
 sky130_fd_sc_hd__and3_1 _12229_ (.A(\cur_mb_mem[172][1] ),
    .B(_06920_),
    .C(_05922_),
    .X(_07274_));
 sky130_fd_sc_hd__and3_2 _12230_ (.A(\cur_mb_mem[26][1] ),
    .B(_05905_),
    .C(_06001_),
    .X(_07275_));
 sky130_fd_sc_hd__a2111o_1 _12231_ (.A1(\cur_mb_mem[42][1] ),
    .A2(_06441_),
    .B1(_07273_),
    .C1(_07274_),
    .D1(_07275_),
    .X(_07276_));
 sky130_fd_sc_hd__buf_8 _12232_ (.A(net253),
    .X(_07277_));
 sky130_fd_sc_hd__and3_1 _12233_ (.A(\cur_mb_mem[93][1] ),
    .B(_07277_),
    .C(_06246_),
    .X(_07278_));
 sky130_fd_sc_hd__buf_12 _12234_ (.A(_06131_),
    .X(_07279_));
 sky130_fd_sc_hd__and3_1 _12235_ (.A(\cur_mb_mem[53][1] ),
    .B(_05056_),
    .C(_07279_),
    .X(_07280_));
 sky130_fd_sc_hd__and3_1 _12236_ (.A(\cur_mb_mem[29][1] ),
    .B(_05945_),
    .C(_05975_),
    .X(_07281_));
 sky130_fd_sc_hd__a2111o_1 _12237_ (.A1(\cur_mb_mem[185][1] ),
    .A2(_06040_),
    .B1(_07278_),
    .C1(_07280_),
    .D1(_07281_),
    .X(_07282_));
 sky130_fd_sc_hd__or4_1 _12238_ (.A(_07268_),
    .B(_07272_),
    .C(_07276_),
    .D(_07282_),
    .X(_07283_));
 sky130_fd_sc_hd__or4_2 _12239_ (.A(_07228_),
    .B(_07246_),
    .C(_07264_),
    .D(_07283_),
    .X(_07284_));
 sky130_fd_sc_hd__or4_4 _12240_ (.A(_07104_),
    .B(_07141_),
    .C(_07211_),
    .D(_07284_),
    .X(_07285_));
 sky130_fd_sc_hd__o22ai_4 _12241_ (.A1(\cur_mb_mem[0][1] ),
    .A2(_05908_),
    .B1(_07028_),
    .B2(_07285_),
    .Y(_07286_));
 sky130_fd_sc_hd__a22o_1 _12242_ (.A1(\cur_mb_mem[223][0] ),
    .A2(_06151_),
    .B1(_06297_),
    .B2(\cur_mb_mem[95][0] ),
    .X(_07287_));
 sky130_fd_sc_hd__a22o_1 _12243_ (.A1(\cur_mb_mem[38][0] ),
    .A2(_06396_),
    .B1(_06075_),
    .B2(\cur_mb_mem[128][0] ),
    .X(_07288_));
 sky130_fd_sc_hd__and3_1 _12244_ (.A(\cur_mb_mem[214][0] ),
    .B(_06186_),
    .C(_05948_),
    .X(_07289_));
 sky130_fd_sc_hd__a31o_4 _12245_ (.A1(\cur_mb_mem[221][0] ),
    .A2(_05946_),
    .A3(_05942_),
    .B1(_07289_),
    .X(_07290_));
 sky130_fd_sc_hd__a211o_1 _12246_ (.A1(\cur_mb_mem[159][0] ),
    .A2(_06174_),
    .B1(_07288_),
    .C1(_07290_),
    .X(_07291_));
 sky130_fd_sc_hd__a221o_1 _12247_ (.A1(\cur_mb_mem[101][0] ),
    .A2(_06269_),
    .B1(_06242_),
    .B2(\cur_mb_mem[22][0] ),
    .C1(_07291_),
    .X(_07292_));
 sky130_fd_sc_hd__a32o_1 _12248_ (.A1(\cur_mb_mem[160][0] ),
    .A2(_06426_),
    .A3(_05973_),
    .B1(_06489_),
    .B2(\cur_mb_mem[25][0] ),
    .X(_07293_));
 sky130_fd_sc_hd__a32o_4 _12249_ (.A1(\cur_mb_mem[148][0] ),
    .A2(_06134_),
    .A3(_05979_),
    .B1(_06322_),
    .B2(\cur_mb_mem[108][0] ),
    .X(_07294_));
 sky130_fd_sc_hd__a221o_1 _12250_ (.A1(\cur_mb_mem[12][0] ),
    .A2(_05928_),
    .B1(_06193_),
    .B2(\cur_mb_mem[166][0] ),
    .C1(_07294_),
    .X(_07295_));
 sky130_fd_sc_hd__a32o_1 _12251_ (.A1(\cur_mb_mem[20][0] ),
    .A2(_06223_),
    .A3(_05976_),
    .B1(_06017_),
    .B2(\cur_mb_mem[28][0] ),
    .X(_07296_));
 sky130_fd_sc_hd__a32o_4 _12252_ (.A1(\cur_mb_mem[219][0] ),
    .A2(_05919_),
    .A3(_05948_),
    .B1(_06040_),
    .B2(\cur_mb_mem[185][0] ),
    .X(_07297_));
 sky130_fd_sc_hd__a22o_1 _12253_ (.A1(\cur_mb_mem[46][0] ),
    .A2(_06107_),
    .B1(_05966_),
    .B2(\cur_mb_mem[129][0] ),
    .X(_07298_));
 sky130_fd_sc_hd__a22o_1 _12254_ (.A1(\cur_mb_mem[45][0] ),
    .A2(_06491_),
    .B1(_06316_),
    .B2(\cur_mb_mem[176][0] ),
    .X(_07299_));
 sky130_fd_sc_hd__a32o_1 _12255_ (.A1(\cur_mb_mem[201][0] ),
    .A2(_05911_),
    .A3(_06092_),
    .B1(_06217_),
    .B2(\cur_mb_mem[180][0] ),
    .X(_07300_));
 sky130_fd_sc_hd__or4_1 _12256_ (.A(_07297_),
    .B(_07298_),
    .C(_07299_),
    .D(_07300_),
    .X(_07301_));
 sky130_fd_sc_hd__or4_1 _12257_ (.A(_07293_),
    .B(_07295_),
    .C(_07296_),
    .D(_07301_),
    .X(_07302_));
 sky130_fd_sc_hd__a2111o_2 _12258_ (.A1(\cur_mb_mem[31][0] ),
    .A2(_06178_),
    .B1(_07287_),
    .C1(_07292_),
    .D1(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__and3_1 _12259_ (.A(\cur_mb_mem[170][0] ),
    .B(_05931_),
    .C(_06758_),
    .X(_07304_));
 sky130_fd_sc_hd__and3_1 _12260_ (.A(\cur_mb_mem[81][0] ),
    .B(_06931_),
    .C(_06353_),
    .X(_07305_));
 sky130_fd_sc_hd__and3_1 _12261_ (.A(\cur_mb_mem[105][0] ),
    .B(_06903_),
    .C(_06268_),
    .X(_07306_));
 sky130_fd_sc_hd__a2111o_2 _12262_ (.A1(\cur_mb_mem[36][0] ),
    .A2(_06360_),
    .B1(_07304_),
    .C1(_07305_),
    .D1(_07306_),
    .X(_07307_));
 sky130_fd_sc_hd__and3_1 _12263_ (.A(\cur_mb_mem[89][0] ),
    .B(_06327_),
    .C(_06378_),
    .X(_07308_));
 sky130_fd_sc_hd__and3_1 _12264_ (.A(\cur_mb_mem[27][0] ),
    .B(_06474_),
    .C(_06235_),
    .X(_07309_));
 sky130_fd_sc_hd__and3_1 _12265_ (.A(\cur_mb_mem[194][0] ),
    .B(_06080_),
    .C(_06082_),
    .X(_07310_));
 sky130_fd_sc_hd__a2111o_1 _12266_ (.A1(\cur_mb_mem[141][0] ),
    .A2(_06250_),
    .B1(_07308_),
    .C1(_07309_),
    .D1(_07310_),
    .X(_07311_));
 sky130_fd_sc_hd__and3_1 _12267_ (.A(\cur_mb_mem[122][0] ),
    .B(_06115_),
    .C(_06051_),
    .X(_07312_));
 sky130_fd_sc_hd__and3_1 _12268_ (.A(\cur_mb_mem[125][0] ),
    .B(_06762_),
    .C(_06138_),
    .X(_07313_));
 sky130_fd_sc_hd__and3_1 _12269_ (.A(\cur_mb_mem[222][0] ),
    .B(_06150_),
    .C(_06000_),
    .X(_07314_));
 sky130_fd_sc_hd__a2111o_2 _12270_ (.A1(\cur_mb_mem[10][0] ),
    .A2(_06408_),
    .B1(_07312_),
    .C1(_07313_),
    .D1(_07314_),
    .X(_07315_));
 sky130_fd_sc_hd__and3_1 _12271_ (.A(\cur_mb_mem[217][0] ),
    .B(_06723_),
    .C(_06814_),
    .X(_07316_));
 sky130_fd_sc_hd__and3_1 _12272_ (.A(\cur_mb_mem[154][0] ),
    .B(_06960_),
    .C(_06747_),
    .X(_07317_));
 sky130_fd_sc_hd__and3_1 _12273_ (.A(\cur_mb_mem[124][0] ),
    .B(_05902_),
    .C(_07253_),
    .X(_07318_));
 sky130_fd_sc_hd__a2111o_2 _12274_ (.A1(\cur_mb_mem[190][0] ),
    .A2(_06480_),
    .B1(_07316_),
    .C1(_07317_),
    .D1(_07318_),
    .X(_07319_));
 sky130_fd_sc_hd__or4_1 _12275_ (.A(_07307_),
    .B(_07311_),
    .C(_07315_),
    .D(_07319_),
    .X(_07320_));
 sky130_fd_sc_hd__and3_1 _12276_ (.A(\cur_mb_mem[57][0] ),
    .B(_06350_),
    .C(_06327_),
    .X(_07321_));
 sky130_fd_sc_hd__and3_1 _12277_ (.A(\cur_mb_mem[86][0] ),
    .B(_05914_),
    .C(_06204_),
    .X(_07322_));
 sky130_fd_sc_hd__and3_1 _12278_ (.A(\cur_mb_mem[136][0] ),
    .B(_05982_),
    .C(_06146_),
    .X(_07323_));
 sky130_fd_sc_hd__a2111o_1 _12279_ (.A1(\cur_mb_mem[4][0] ),
    .A2(_06162_),
    .B1(_07321_),
    .C1(_07322_),
    .D1(_07323_),
    .X(_07324_));
 sky130_fd_sc_hd__and3_4 _12280_ (.A(\cur_mb_mem[192][0] ),
    .B(_06456_),
    .C(_06009_),
    .X(_07325_));
 sky130_fd_sc_hd__and3_1 _12281_ (.A(\cur_mb_mem[77][0] ),
    .B(_06490_),
    .C(_06809_),
    .X(_07326_));
 sky130_fd_sc_hd__and3_2 _12282_ (.A(\cur_mb_mem[58][0] ),
    .B(_06198_),
    .C(_06960_),
    .X(_07327_));
 sky130_fd_sc_hd__a2111o_1 _12283_ (.A1(\cur_mb_mem[132][0] ),
    .A2(net220),
    .B1(_07325_),
    .C1(_07326_),
    .D1(_07327_),
    .X(_07328_));
 sky130_fd_sc_hd__and3_1 _12284_ (.A(\cur_mb_mem[69][0] ),
    .B(_06233_),
    .C(_06812_),
    .X(_07329_));
 sky130_fd_sc_hd__and3_4 _12285_ (.A(\cur_mb_mem[51][0] ),
    .B(_06240_),
    .C(_06770_),
    .X(_07330_));
 sky130_fd_sc_hd__and3_1 _12286_ (.A(\cur_mb_mem[64][0] ),
    .B(_06057_),
    .C(_06748_),
    .X(_07331_));
 sky130_fd_sc_hd__a2111o_1 _12287_ (.A1(\cur_mb_mem[29][0] ),
    .A2(_06404_),
    .B1(_07329_),
    .C1(_07330_),
    .D1(_07331_),
    .X(_07332_));
 sky130_fd_sc_hd__and3_1 _12288_ (.A(\cur_mb_mem[70][0] ),
    .B(_06199_),
    .C(_06809_),
    .X(_07333_));
 sky130_fd_sc_hd__and3_1 _12289_ (.A(\cur_mb_mem[65][0] ),
    .B(_06057_),
    .C(_06912_),
    .X(_07334_));
 sky130_fd_sc_hd__and3_1 _12290_ (.A(\cur_mb_mem[78][0] ),
    .B(_06023_),
    .C(_07084_),
    .X(_07335_));
 sky130_fd_sc_hd__a2111o_1 _12291_ (.A1(\cur_mb_mem[19][0] ),
    .A2(_06282_),
    .B1(_07333_),
    .C1(_07334_),
    .D1(_07335_),
    .X(_07336_));
 sky130_fd_sc_hd__or4_4 _12292_ (.A(_07324_),
    .B(_07328_),
    .C(_07332_),
    .D(_07336_),
    .X(_07337_));
 sky130_fd_sc_hd__and3_1 _12293_ (.A(\cur_mb_mem[85][0] ),
    .B(_06931_),
    .C(_06812_),
    .X(_07338_));
 sky130_fd_sc_hd__and3_1 _12294_ (.A(\cur_mb_mem[171][0] ),
    .B(_06474_),
    .C(_06755_),
    .X(_07339_));
 sky130_fd_sc_hd__and3_1 _12295_ (.A(\cur_mb_mem[1][0] ),
    .B(_07096_),
    .C(_06251_),
    .X(_07340_));
 sky130_fd_sc_hd__a2111o_2 _12296_ (.A1(\cur_mb_mem[100][0] ),
    .A2(_06028_),
    .B1(_07338_),
    .C1(_07339_),
    .D1(_07340_),
    .X(_07341_));
 sky130_fd_sc_hd__and3_1 _12297_ (.A(\cur_mb_mem[116][0] ),
    .B(net260),
    .C(_06731_),
    .X(_07342_));
 sky130_fd_sc_hd__and3_1 _12298_ (.A(\cur_mb_mem[202][0] ),
    .B(_05904_),
    .C(_06789_),
    .X(_07343_));
 sky130_fd_sc_hd__and3_1 _12299_ (.A(\cur_mb_mem[252][0] ),
    .B(_06032_),
    .C(_05901_),
    .X(_07344_));
 sky130_fd_sc_hd__and3_1 _12300_ (.A(\cur_mb_mem[13][0] ),
    .B(_06365_),
    .C(_06033_),
    .X(_07345_));
 sky130_fd_sc_hd__or4_1 _12301_ (.A(_07342_),
    .B(_07343_),
    .C(_07344_),
    .D(_07345_),
    .X(_07346_));
 sky130_fd_sc_hd__and3_1 _12302_ (.A(\cur_mb_mem[181][0] ),
    .B(_06760_),
    .C(_06147_),
    .X(_07347_));
 sky130_fd_sc_hd__and3_1 _12303_ (.A(\cur_mb_mem[209][0] ),
    .B(_06814_),
    .C(_06912_),
    .X(_07348_));
 sky130_fd_sc_hd__and3_1 _12304_ (.A(\cur_mb_mem[200][0] ),
    .B(_06832_),
    .C(_06997_),
    .X(_07349_));
 sky130_fd_sc_hd__a2111o_2 _12305_ (.A1(\cur_mb_mem[14][0] ),
    .A2(_06367_),
    .B1(_07347_),
    .C1(_07348_),
    .D1(_07349_),
    .X(_07350_));
 sky130_fd_sc_hd__and3_1 _12306_ (.A(\cur_mb_mem[165][0] ),
    .B(_06192_),
    .C(_06794_),
    .X(_07351_));
 sky130_fd_sc_hd__and3_1 _12307_ (.A(\cur_mb_mem[126][0] ),
    .B(_07078_),
    .C(_06000_),
    .X(_07352_));
 sky130_fd_sc_hd__and3_1 _12308_ (.A(\cur_mb_mem[73][0] ),
    .B(_06834_),
    .C(_06023_),
    .X(_07353_));
 sky130_fd_sc_hd__a2111o_2 _12309_ (.A1(\cur_mb_mem[67][0] ),
    .A2(_06429_),
    .B1(_07351_),
    .C1(_07352_),
    .D1(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__or4_1 _12310_ (.A(_07341_),
    .B(_07346_),
    .C(_07350_),
    .D(_07354_),
    .X(_07355_));
 sky130_fd_sc_hd__and3_1 _12311_ (.A(\cur_mb_mem[9][0] ),
    .B(_06707_),
    .C(_06723_),
    .X(_07356_));
 sky130_fd_sc_hd__and3_1 _12312_ (.A(\cur_mb_mem[145][0] ),
    .B(_06747_),
    .C(_06912_),
    .X(_07357_));
 sky130_fd_sc_hd__and3_1 _12313_ (.A(\cur_mb_mem[158][0] ),
    .B(_07100_),
    .C(_07084_),
    .X(_07358_));
 sky130_fd_sc_hd__a2111o_2 _12314_ (.A1(\cur_mb_mem[203][0] ),
    .A2(_06325_),
    .B1(_07356_),
    .C1(_07357_),
    .D1(_07358_),
    .X(_07359_));
 sky130_fd_sc_hd__and3_1 _12315_ (.A(\cur_mb_mem[34][0] ),
    .B(_06080_),
    .C(_06952_),
    .X(_07360_));
 sky130_fd_sc_hd__and3_1 _12316_ (.A(\cur_mb_mem[186][0] ),
    .B(_06960_),
    .C(_06877_),
    .X(_07361_));
 sky130_fd_sc_hd__and3_1 _12317_ (.A(\cur_mb_mem[16][0] ),
    .B(_06315_),
    .C(_06001_),
    .X(_07362_));
 sky130_fd_sc_hd__a2111o_2 _12318_ (.A1(\cur_mb_mem[11][0] ),
    .A2(_06301_),
    .B1(_07360_),
    .C1(_07361_),
    .D1(_07362_),
    .X(_07363_));
 sky130_fd_sc_hd__and3_1 _12319_ (.A(\cur_mb_mem[35][0] ),
    .B(_06770_),
    .C(_06952_),
    .X(_07364_));
 sky130_fd_sc_hd__and3_1 _12320_ (.A(\cur_mb_mem[54][0] ),
    .B(_07235_),
    .C(_06191_),
    .X(_07365_));
 sky130_fd_sc_hd__and3_2 _12321_ (.A(\cur_mb_mem[204][0] ),
    .B(_06920_),
    .C(_06091_),
    .X(_07366_));
 sky130_fd_sc_hd__a2111o_4 _12322_ (.A1(\cur_mb_mem[131][0] ),
    .A2(_06383_),
    .B1(_07364_),
    .C1(_07365_),
    .D1(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__and3_2 _12323_ (.A(\cur_mb_mem[244][0] ),
    .B(_07137_),
    .C(_06215_),
    .X(_07368_));
 sky130_fd_sc_hd__and3_1 _12324_ (.A(\cur_mb_mem[3][0] ),
    .B(_07096_),
    .C(_06086_),
    .X(_07369_));
 sky130_fd_sc_hd__and3_1 _12325_ (.A(\cur_mb_mem[113][0] ),
    .B(_07021_),
    .C(_05993_),
    .X(_07370_));
 sky130_fd_sc_hd__a2111o_1 _12326_ (.A1(\cur_mb_mem[155][0] ),
    .A2(_06402_),
    .B1(_07368_),
    .C1(_07369_),
    .D1(_07370_),
    .X(_07371_));
 sky130_fd_sc_hd__or4_1 _12327_ (.A(_07359_),
    .B(_07363_),
    .C(_07367_),
    .D(_07371_),
    .X(_07372_));
 sky130_fd_sc_hd__or4_4 _12328_ (.A(_07320_),
    .B(_07337_),
    .C(_07355_),
    .D(_07372_),
    .X(_07373_));
 sky130_fd_sc_hd__a32o_1 _12329_ (.A1(\cur_mb_mem[247][0] ),
    .A2(_04430_),
    .A3(_06096_),
    .B1(_06248_),
    .B2(\cur_mb_mem[237][0] ),
    .X(_07374_));
 sky130_fd_sc_hd__a32o_1 _12330_ (.A1(\cur_mb_mem[175][0] ),
    .A2(_04423_),
    .A3(_06137_),
    .B1(_06447_),
    .B2(\cur_mb_mem[215][0] ),
    .X(_07375_));
 sky130_fd_sc_hd__a2111o_2 _12331_ (.A1(\cur_mb_mem[127][0] ),
    .A2(_06101_),
    .B1(_07374_),
    .C1(_07375_),
    .D1(_06185_),
    .X(_07376_));
 sky130_fd_sc_hd__a22o_1 _12332_ (.A1(\cur_mb_mem[242][0] ),
    .A2(_06335_),
    .B1(_06195_),
    .B2(\cur_mb_mem[164][0] ),
    .X(_07377_));
 sky130_fd_sc_hd__a221o_1 _12333_ (.A1(\cur_mb_mem[216][0] ),
    .A2(_06317_),
    .B1(_06433_),
    .B2(\cur_mb_mem[144][0] ),
    .C1(_07377_),
    .X(_07378_));
 sky130_fd_sc_hd__a22o_1 _12334_ (.A1(\cur_mb_mem[226][0] ),
    .A2(_06256_),
    .B1(_06180_),
    .B2(\cur_mb_mem[231][0] ),
    .X(_07379_));
 sky130_fd_sc_hd__a32o_1 _12335_ (.A1(\cur_mb_mem[235][0] ),
    .A2(_06261_),
    .A3(_06224_),
    .B1(_06344_),
    .B2(\cur_mb_mem[37][0] ),
    .X(_07380_));
 sky130_fd_sc_hd__and3_1 _12336_ (.A(\cur_mb_mem[15][0] ),
    .B(_06466_),
    .C(_06202_),
    .X(_07381_));
 sky130_fd_sc_hd__and3_1 _12337_ (.A(\cur_mb_mem[232][0] ),
    .B(_05982_),
    .C(_06247_),
    .X(_07382_));
 sky130_fd_sc_hd__and3_1 _12338_ (.A(\cur_mb_mem[234][0] ),
    .B(_05905_),
    .C(_06918_),
    .X(_07383_));
 sky130_fd_sc_hd__a2111o_1 _12339_ (.A1(\cur_mb_mem[134][0] ),
    .A2(_06211_),
    .B1(_07381_),
    .C1(_07382_),
    .D1(_07383_),
    .X(_07384_));
 sky130_fd_sc_hd__and3_1 _12340_ (.A(\cur_mb_mem[246][0] ),
    .B(_06902_),
    .C(_06199_),
    .X(_07385_));
 sky130_fd_sc_hd__and3_1 _12341_ (.A(\cur_mb_mem[227][0] ),
    .B(_06980_),
    .C(_06918_),
    .X(_07386_));
 sky130_fd_sc_hd__and3_1 _12342_ (.A(\cur_mb_mem[184][0] ),
    .B(_06774_),
    .C(_06216_),
    .X(_07387_));
 sky130_fd_sc_hd__a2111o_1 _12343_ (.A1(\cur_mb_mem[177][0] ),
    .A2(_06020_),
    .B1(_07385_),
    .C1(_07386_),
    .D1(_07387_),
    .X(_07388_));
 sky130_fd_sc_hd__or4_2 _12344_ (.A(_07379_),
    .B(_07380_),
    .C(_07384_),
    .D(_07388_),
    .X(_07389_));
 sky130_fd_sc_hd__and3_1 _12345_ (.A(\cur_mb_mem[172][0] ),
    .B(_06754_),
    .C(_06755_),
    .X(_07390_));
 sky130_fd_sc_hd__and3_1 _12346_ (.A(\cur_mb_mem[43][0] ),
    .B(_06387_),
    .C(_06087_),
    .X(_07391_));
 sky130_fd_sc_hd__and3_1 _12347_ (.A(\cur_mb_mem[88][0] ),
    .B(_06774_),
    .C(_07277_),
    .X(_07392_));
 sky130_fd_sc_hd__a2111o_1 _12348_ (.A1(\cur_mb_mem[61][0] ),
    .A2(_06359_),
    .B1(_07390_),
    .C1(_07391_),
    .D1(_07392_),
    .X(_07393_));
 sky130_fd_sc_hd__and3_2 _12349_ (.A(\cur_mb_mem[245][0] ),
    .B(_06916_),
    .C(_06208_),
    .X(_07394_));
 sky130_fd_sc_hd__and3_1 _12350_ (.A(\cur_mb_mem[112][0] ),
    .B(_07078_),
    .C(_06748_),
    .X(_07395_));
 sky130_fd_sc_hd__and3_1 _12351_ (.A(\cur_mb_mem[72][0] ),
    .B(_06774_),
    .C(_06023_),
    .X(_07396_));
 sky130_fd_sc_hd__a2111o_1 _12352_ (.A1(\cur_mb_mem[138][0] ),
    .A2(_05934_),
    .B1(_07394_),
    .C1(_07395_),
    .D1(_07396_),
    .X(_07397_));
 sky130_fd_sc_hd__and3_1 _12353_ (.A(\cur_mb_mem[133][0] ),
    .B(_06859_),
    .C(_06794_),
    .X(_07398_));
 sky130_fd_sc_hd__and3_1 _12354_ (.A(\cur_mb_mem[117][0] ),
    .B(_07078_),
    .C(_06153_),
    .X(_07399_));
 sky130_fd_sc_hd__and3_1 _12355_ (.A(\cur_mb_mem[120][0] ),
    .B(_06774_),
    .C(_07253_),
    .X(_07400_));
 sky130_fd_sc_hd__a2111o_1 _12356_ (.A1(\cur_mb_mem[97][0] ),
    .A2(_06077_),
    .B1(_07398_),
    .C1(_07399_),
    .D1(_07400_),
    .X(_07401_));
 sky130_fd_sc_hd__and3_1 _12357_ (.A(\cur_mb_mem[196][0] ),
    .B(_06026_),
    .C(_06324_),
    .X(_07402_));
 sky130_fd_sc_hd__and3_1 _12358_ (.A(\cur_mb_mem[198][0] ),
    .B(_06210_),
    .C(_06456_),
    .X(_07403_));
 sky130_fd_sc_hd__and3_1 _12359_ (.A(\cur_mb_mem[208][0] ),
    .B(_06348_),
    .C(_06009_),
    .X(_07404_));
 sky130_fd_sc_hd__and3_4 _12360_ (.A(\cur_mb_mem[75][0] ),
    .B(_06474_),
    .C(_06809_),
    .X(_07405_));
 sky130_fd_sc_hd__or4_4 _12361_ (.A(_07402_),
    .B(_07403_),
    .C(_07404_),
    .D(_07405_),
    .X(_07406_));
 sky130_fd_sc_hd__or4_4 _12362_ (.A(_07393_),
    .B(_07397_),
    .C(_07401_),
    .D(_07406_),
    .X(_07407_));
 sky130_fd_sc_hd__or4_1 _12363_ (.A(_07376_),
    .B(_07378_),
    .C(_07389_),
    .D(_07407_),
    .X(_07408_));
 sky130_fd_sc_hd__and3_1 _12364_ (.A(\cur_mb_mem[169][0] ),
    .B(_06327_),
    .C(_06825_),
    .X(_07409_));
 sky130_fd_sc_hd__and3_1 _12365_ (.A(\cur_mb_mem[168][0] ),
    .B(_06478_),
    .C(_06825_),
    .X(_07410_));
 sky130_fd_sc_hd__and3_1 _12366_ (.A(\cur_mb_mem[33][0] ),
    .B(_06087_),
    .C(_06251_),
    .X(_07411_));
 sky130_fd_sc_hd__a2111o_1 _12367_ (.A1(\cur_mb_mem[42][0] ),
    .A2(_06441_),
    .B1(_07409_),
    .C1(_07410_),
    .D1(_07411_),
    .X(_07412_));
 sky130_fd_sc_hd__and3_1 _12368_ (.A(\cur_mb_mem[102][0] ),
    .B(_05984_),
    .C(_06140_),
    .X(_07413_));
 sky130_fd_sc_hd__and3_1 _12369_ (.A(\cur_mb_mem[193][0] ),
    .B(_06352_),
    .C(_06841_),
    .X(_07414_));
 sky130_fd_sc_hd__and3_1 _12370_ (.A(\cur_mb_mem[96][0] ),
    .B(_06268_),
    .C(_06748_),
    .X(_07415_));
 sky130_fd_sc_hd__a2111o_1 _12371_ (.A1(\cur_mb_mem[74][0] ),
    .A2(_06417_),
    .B1(_07413_),
    .C1(_07414_),
    .D1(_07415_),
    .X(_07416_));
 sky130_fd_sc_hd__and3_2 _12372_ (.A(\cur_mb_mem[218][0] ),
    .B(_05957_),
    .C(_06814_),
    .X(_07417_));
 sky130_fd_sc_hd__and3_1 _12373_ (.A(\cur_mb_mem[137][0] ),
    .B(_06903_),
    .C(_06146_),
    .X(_07418_));
 sky130_fd_sc_hd__and3_1 _12374_ (.A(\cur_mb_mem[179][0] ),
    .B(_06980_),
    .C(_06877_),
    .X(_07419_));
 sky130_fd_sc_hd__a2111o_1 _12375_ (.A1(\cur_mb_mem[152][0] ),
    .A2(_06394_),
    .B1(_07417_),
    .C1(_07418_),
    .D1(_07419_),
    .X(_07420_));
 sky130_fd_sc_hd__and3_1 _12376_ (.A(\cur_mb_mem[109][0] ),
    .B(_06268_),
    .C(_06056_),
    .X(_07421_));
 sky130_fd_sc_hd__and3_1 _12377_ (.A(\cur_mb_mem[84][0] ),
    .B(_06215_),
    .C(_06895_),
    .X(_07422_));
 sky130_fd_sc_hd__and3_1 _12378_ (.A(\cur_mb_mem[251][0] ),
    .B(_07137_),
    .C(_05918_),
    .X(_07423_));
 sky130_fd_sc_hd__a2111o_1 _12379_ (.A1(\cur_mb_mem[110][0] ),
    .A2(_06047_),
    .B1(_07421_),
    .C1(_07422_),
    .D1(_07423_),
    .X(_07424_));
 sky130_fd_sc_hd__or4_2 _12380_ (.A(_07412_),
    .B(_07416_),
    .C(_07420_),
    .D(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__and3_1 _12381_ (.A(\cur_mb_mem[80][0] ),
    .B(_06931_),
    .C(_06815_),
    .X(_07426_));
 sky130_fd_sc_hd__and3_1 _12382_ (.A(\cur_mb_mem[17][0] ),
    .B(_06841_),
    .C(_06235_),
    .X(_07427_));
 sky130_fd_sc_hd__and3_1 _12383_ (.A(\cur_mb_mem[62][0] ),
    .B(_06198_),
    .C(_06000_),
    .X(_07428_));
 sky130_fd_sc_hd__a2111o_2 _12384_ (.A1(\cur_mb_mem[24][0] ),
    .A2(_06285_),
    .B1(_07426_),
    .C1(_07427_),
    .D1(_07428_),
    .X(_07429_));
 sky130_fd_sc_hd__and3_1 _12385_ (.A(\cur_mb_mem[130][0] ),
    .B(_06254_),
    .C(_06842_),
    .X(_07430_));
 sky130_fd_sc_hd__and3_2 _12386_ (.A(\cur_mb_mem[197][0] ),
    .B(_06352_),
    .C(_06208_),
    .X(_07431_));
 sky130_fd_sc_hd__and3_1 _12387_ (.A(\cur_mb_mem[92][0] ),
    .B(_06937_),
    .C(_06895_),
    .X(_07432_));
 sky130_fd_sc_hd__a2111o_1 _12388_ (.A1(\cur_mb_mem[161][0] ),
    .A2(_06334_),
    .B1(_07430_),
    .C1(_07431_),
    .D1(_07432_),
    .X(_07433_));
 sky130_fd_sc_hd__and3_2 _12389_ (.A(\cur_mb_mem[106][0] ),
    .B(_05957_),
    .C(_05984_),
    .X(_07434_));
 sky130_fd_sc_hd__and3_1 _12390_ (.A(\cur_mb_mem[188][0] ),
    .B(_06754_),
    .C(_06830_),
    .X(_07435_));
 sky130_fd_sc_hd__and3_1 _12391_ (.A(\cur_mb_mem[82][0] ),
    .B(_06380_),
    .C(_06895_),
    .X(_07436_));
 sky130_fd_sc_hd__a2111o_1 _12392_ (.A1(\cur_mb_mem[44][0] ),
    .A2(_06399_),
    .B1(_07434_),
    .C1(_07435_),
    .D1(_07436_),
    .X(_07437_));
 sky130_fd_sc_hd__and3_1 _12393_ (.A(\cur_mb_mem[254][0] ),
    .B(_06902_),
    .C(_06000_),
    .X(_07438_));
 sky130_fd_sc_hd__and3_1 _12394_ (.A(\cur_mb_mem[150][0] ),
    .B(_06191_),
    .C(_06152_),
    .X(_07439_));
 sky130_fd_sc_hd__and3_1 _12395_ (.A(\cur_mb_mem[212][0] ),
    .B(_05890_),
    .C(_05947_),
    .X(_07440_));
 sky130_fd_sc_hd__a2111o_4 _12396_ (.A1(\cur_mb_mem[253][0] ),
    .A2(_06034_),
    .B1(_07438_),
    .C1(_07439_),
    .D1(_07440_),
    .X(_07441_));
 sky130_fd_sc_hd__or4_2 _12397_ (.A(_07429_),
    .B(_07433_),
    .C(_07437_),
    .D(_07441_),
    .X(_07442_));
 sky130_fd_sc_hd__and3_1 _12398_ (.A(\cur_mb_mem[93][0] ),
    .B(_05913_),
    .C(_06033_),
    .X(_07443_));
 sky130_fd_sc_hd__and3_1 _12399_ (.A(\cur_mb_mem[220][0] ),
    .B(_06321_),
    .C(_06802_),
    .X(_07444_));
 sky130_fd_sc_hd__and3_1 _12400_ (.A(\cur_mb_mem[174][0] ),
    .B(_05953_),
    .C(_06333_),
    .X(_07445_));
 sky130_fd_sc_hd__and3_1 _12401_ (.A(\cur_mb_mem[206][0] ),
    .B(_06366_),
    .C(_06986_),
    .X(_07446_));
 sky130_fd_sc_hd__or4_1 _12402_ (.A(_07443_),
    .B(_07444_),
    .C(_07445_),
    .D(_07446_),
    .X(_07447_));
 sky130_fd_sc_hd__and3_4 _12403_ (.A(\cur_mb_mem[32][0] ),
    .B(_06343_),
    .C(_05970_),
    .X(_07448_));
 sky130_fd_sc_hd__and3_1 _12404_ (.A(\cur_mb_mem[8][0] ),
    .B(_06707_),
    .C(_05982_),
    .X(_07449_));
 sky130_fd_sc_hd__and3_1 _12405_ (.A(\cur_mb_mem[156][0] ),
    .B(_05902_),
    .C(_06152_),
    .X(_07450_));
 sky130_fd_sc_hd__a2111o_1 _12406_ (.A1(\cur_mb_mem[211][0] ),
    .A2(_06349_),
    .B1(_07448_),
    .C1(_07449_),
    .D1(_07450_),
    .X(_07451_));
 sky130_fd_sc_hd__and3_1 _12407_ (.A(\cur_mb_mem[157][0] ),
    .B(_06762_),
    .C(_06747_),
    .X(_07452_));
 sky130_fd_sc_hd__and3_1 _12408_ (.A(\cur_mb_mem[21][0] ),
    .B(_06235_),
    .C(_06794_),
    .X(_07453_));
 sky130_fd_sc_hd__and3_1 _12409_ (.A(\cur_mb_mem[249][0] ),
    .B(_07137_),
    .C(_06834_),
    .X(_07454_));
 sky130_fd_sc_hd__a2111o_1 _12410_ (.A1(\cur_mb_mem[250][0] ),
    .A2(_06443_),
    .B1(_07452_),
    .C1(_07453_),
    .D1(_07454_),
    .X(_07455_));
 sky130_fd_sc_hd__and3_1 _12411_ (.A(\cur_mb_mem[213][0] ),
    .B(_06150_),
    .C(_06153_),
    .X(_07456_));
 sky130_fd_sc_hd__and3_1 _12412_ (.A(\cur_mb_mem[149][0] ),
    .B(_07100_),
    .C(_07279_),
    .X(_07457_));
 sky130_fd_sc_hd__and3_1 _12413_ (.A(\cur_mb_mem[107][0] ),
    .B(_05918_),
    .C(_06413_),
    .X(_07458_));
 sky130_fd_sc_hd__a2111o_1 _12414_ (.A1(\cur_mb_mem[6][0] ),
    .A2(_06203_),
    .B1(_07456_),
    .C1(_07457_),
    .D1(_07458_),
    .X(_07459_));
 sky130_fd_sc_hd__or4_4 _12415_ (.A(_07447_),
    .B(_07451_),
    .C(_07455_),
    .D(_07459_),
    .X(_07460_));
 sky130_fd_sc_hd__and3_1 _12416_ (.A(\cur_mb_mem[243][0] ),
    .B(_06916_),
    .C(_06770_),
    .X(_07461_));
 sky130_fd_sc_hd__and3_1 _12417_ (.A(\cur_mb_mem[229][0] ),
    .B(_06153_),
    .C(_06918_),
    .X(_07462_));
 sky130_fd_sc_hd__and3_1 _12418_ (.A(\cur_mb_mem[60][0] ),
    .B(_05056_),
    .C(_06920_),
    .X(_07463_));
 sky130_fd_sc_hd__a2111o_1 _12419_ (.A1(\cur_mb_mem[53][0] ),
    .A2(_06221_),
    .B1(_07461_),
    .C1(_07462_),
    .D1(_07463_),
    .X(_07464_));
 sky130_fd_sc_hd__and3_1 _12420_ (.A(\cur_mb_mem[207][0] ),
    .B(_06149_),
    .C(_06967_),
    .X(_07465_));
 sky130_fd_sc_hd__and3_1 _12421_ (.A(\cur_mb_mem[236][0] ),
    .B(_05902_),
    .C(_06918_),
    .X(_07466_));
 sky130_fd_sc_hd__and3_1 _12422_ (.A(\cur_mb_mem[167][0] ),
    .B(_05922_),
    .C(_06096_),
    .X(_07467_));
 sky130_fd_sc_hd__a2111o_1 _12423_ (.A1(\cur_mb_mem[79][0] ),
    .A2(_06122_),
    .B1(_07465_),
    .C1(_07466_),
    .D1(_07467_),
    .X(_07468_));
 sky130_fd_sc_hd__and3_1 _12424_ (.A(\cur_mb_mem[48][0] ),
    .B(_06198_),
    .C(_06748_),
    .X(_07469_));
 sky130_fd_sc_hd__and3_1 _12425_ (.A(\cur_mb_mem[241][0] ),
    .B(_07137_),
    .C(_06251_),
    .X(_07470_));
 sky130_fd_sc_hd__and3_1 _12426_ (.A(\cur_mb_mem[41][0] ),
    .B(_05893_),
    .C(_06044_),
    .X(_07471_));
 sky130_fd_sc_hd__a2111o_1 _12427_ (.A1(\cur_mb_mem[182][0] ),
    .A2(_06205_),
    .B1(_07469_),
    .C1(_07470_),
    .D1(_07471_),
    .X(_07472_));
 sky130_fd_sc_hd__and3_4 _12428_ (.A(\cur_mb_mem[26][0] ),
    .B(_05931_),
    .C(_06475_),
    .X(_07473_));
 sky130_fd_sc_hd__and3_1 _12429_ (.A(\cur_mb_mem[240][0] ),
    .B(_06158_),
    .C(_06009_),
    .X(_07474_));
 sky130_fd_sc_hd__and3_1 _12430_ (.A(\cur_mb_mem[183][0] ),
    .B(_06019_),
    .C(_06179_),
    .X(_07475_));
 sky130_fd_sc_hd__and3_1 _12431_ (.A(\cur_mb_mem[23][0] ),
    .B(_06708_),
    .C(_06235_),
    .X(_07476_));
 sky130_fd_sc_hd__or4_1 _12432_ (.A(_07473_),
    .B(_07474_),
    .C(_07475_),
    .D(_07476_),
    .X(_07477_));
 sky130_fd_sc_hd__or4_4 _12433_ (.A(_07464_),
    .B(_07468_),
    .C(_07472_),
    .D(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__or4_2 _12434_ (.A(_07425_),
    .B(_07442_),
    .C(_07460_),
    .D(_07478_),
    .X(_07479_));
 sky130_fd_sc_hd__and3_1 _12435_ (.A(\cur_mb_mem[63][0] ),
    .B(_06466_),
    .C(_06240_),
    .X(_07480_));
 sky130_fd_sc_hd__and3_1 _12436_ (.A(\cur_mb_mem[224][0] ),
    .B(_06772_),
    .C(_06247_),
    .X(_07481_));
 sky130_fd_sc_hd__and3_1 _12437_ (.A(\cur_mb_mem[191][0] ),
    .B(_04423_),
    .C(_06877_),
    .X(_07482_));
 sky130_fd_sc_hd__a2111o_4 _12438_ (.A1(\cur_mb_mem[255][0] ),
    .A2(_06304_),
    .B1(_07480_),
    .C1(_07481_),
    .D1(_07482_),
    .X(_07483_));
 sky130_fd_sc_hd__and3_1 _12439_ (.A(\cur_mb_mem[111][0] ),
    .B(_06099_),
    .C(_06267_),
    .X(_07484_));
 sky130_fd_sc_hd__and3_1 _12440_ (.A(\cur_mb_mem[71][0] ),
    .B(_06022_),
    .C(_06851_),
    .X(_07485_));
 sky130_fd_sc_hd__and3_1 _12441_ (.A(\cur_mb_mem[103][0] ),
    .B(_06027_),
    .C(_06461_),
    .X(_07486_));
 sky130_fd_sc_hd__and3_1 _12442_ (.A(\cur_mb_mem[47][0] ),
    .B(_06120_),
    .C(_06395_),
    .X(_07487_));
 sky130_fd_sc_hd__or4_4 _12443_ (.A(_07484_),
    .B(_07485_),
    .C(_07486_),
    .D(_07487_),
    .X(_07488_));
 sky130_fd_sc_hd__and3_1 _12444_ (.A(\cur_mb_mem[40][0] ),
    .B(_06832_),
    .C(_06952_),
    .X(_07489_));
 sky130_fd_sc_hd__and3_1 _12445_ (.A(\cur_mb_mem[98][0] ),
    .B(_06908_),
    .C(_06413_),
    .X(_07490_));
 sky130_fd_sc_hd__and3_1 _12446_ (.A(\cur_mb_mem[210][0] ),
    .B(_07099_),
    .C(_05947_),
    .X(_07491_));
 sky130_fd_sc_hd__a2111o_1 _12447_ (.A1(\cur_mb_mem[91][0] ),
    .A2(_06361_),
    .B1(_07489_),
    .C1(_07490_),
    .D1(_07491_),
    .X(_07492_));
 sky130_fd_sc_hd__and3_4 _12448_ (.A(\cur_mb_mem[238][0] ),
    .B(_07084_),
    .C(_06918_),
    .X(_07493_));
 sky130_fd_sc_hd__and3_1 _12449_ (.A(\cur_mb_mem[151][0] ),
    .B(_07100_),
    .C(_06096_),
    .X(_07494_));
 sky130_fd_sc_hd__and3_1 _12450_ (.A(\cur_mb_mem[123][0] ),
    .B(_05918_),
    .C(_07021_),
    .X(_07495_));
 sky130_fd_sc_hd__a2111o_1 _12451_ (.A1(\cur_mb_mem[68][0] ),
    .A2(_06234_),
    .B1(_07493_),
    .C1(_07494_),
    .D1(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__or4_4 _12452_ (.A(_07483_),
    .B(_07488_),
    .C(_07492_),
    .D(_07496_),
    .X(_07497_));
 sky130_fd_sc_hd__and3_2 _12453_ (.A(\cur_mb_mem[146][0] ),
    .B(_06080_),
    .C(_06747_),
    .X(_07498_));
 sky130_fd_sc_hd__and3_1 _12454_ (.A(\cur_mb_mem[199][0] ),
    .B(_06967_),
    .C(_06896_),
    .X(_07499_));
 sky130_fd_sc_hd__and3_1 _12455_ (.A(\cur_mb_mem[87][0] ),
    .B(_07277_),
    .C(_07195_),
    .X(_07500_));
 sky130_fd_sc_hd__a2111o_1 _12456_ (.A1(\cur_mb_mem[135][0] ),
    .A2(_06462_),
    .B1(_07498_),
    .C1(_07499_),
    .D1(_07500_),
    .X(_07501_));
 sky130_fd_sc_hd__and3_1 _12457_ (.A(\cur_mb_mem[76][0] ),
    .B(_06754_),
    .C(_06809_),
    .X(_07502_));
 sky130_fd_sc_hd__and3_4 _12458_ (.A(\cur_mb_mem[114][0] ),
    .B(_06908_),
    .C(_07078_),
    .X(_07503_));
 sky130_fd_sc_hd__and3_1 _12459_ (.A(\cur_mb_mem[49][0] ),
    .B(_07235_),
    .C(_06251_),
    .X(_07504_));
 sky130_fd_sc_hd__a2111o_1 _12460_ (.A1(\cur_mb_mem[225][0] ),
    .A2(_05998_),
    .B1(_07502_),
    .C1(_07503_),
    .D1(_07504_),
    .X(_07505_));
 sky130_fd_sc_hd__and3_1 _12461_ (.A(\cur_mb_mem[7][0] ),
    .B(_06707_),
    .C(_06708_),
    .X(_07506_));
 sky130_fd_sc_hd__and3_1 _12462_ (.A(\cur_mb_mem[119][0] ),
    .B(_07078_),
    .C(_06896_),
    .X(_07507_));
 sky130_fd_sc_hd__and3_1 _12463_ (.A(\cur_mb_mem[233][0] ),
    .B(_05893_),
    .C(_06065_),
    .X(_07508_));
 sky130_fd_sc_hd__a2111o_1 _12464_ (.A1(\cur_mb_mem[248][0] ),
    .A2(_06411_),
    .B1(_07506_),
    .C1(_07507_),
    .D1(_07508_),
    .X(_07509_));
 sky130_fd_sc_hd__and3_1 _12465_ (.A(\cur_mb_mem[55][0] ),
    .B(_07235_),
    .C(_07195_),
    .X(_07510_));
 sky130_fd_sc_hd__and3_1 _12466_ (.A(\cur_mb_mem[143][0] ),
    .B(_04423_),
    .C(_05935_),
    .X(_07511_));
 sky130_fd_sc_hd__and3_1 _12467_ (.A(\cur_mb_mem[228][0] ),
    .B(_05890_),
    .C(_06065_),
    .X(_07512_));
 sky130_fd_sc_hd__a2111o_1 _12468_ (.A1(\cur_mb_mem[39][0] ),
    .A2(_06373_),
    .B1(_07510_),
    .C1(_07511_),
    .D1(_07512_),
    .X(_07513_));
 sky130_fd_sc_hd__or4_2 _12469_ (.A(_07501_),
    .B(_07505_),
    .C(_07509_),
    .D(_07513_),
    .X(_07514_));
 sky130_fd_sc_hd__and3_1 _12470_ (.A(\cur_mb_mem[173][0] ),
    .B(_06056_),
    .C(_06192_),
    .X(_07515_));
 sky130_fd_sc_hd__and3_1 _12471_ (.A(\cur_mb_mem[205][0] ),
    .B(_06056_),
    .C(_06997_),
    .X(_07516_));
 sky130_fd_sc_hd__and3_1 _12472_ (.A(\cur_mb_mem[139][0] ),
    .B(_06942_),
    .C(_05935_),
    .X(_07517_));
 sky130_fd_sc_hd__a2111o_2 _12473_ (.A1(\cur_mb_mem[142][0] ),
    .A2(_06487_),
    .B1(_07515_),
    .C1(_07516_),
    .D1(_07517_),
    .X(_07518_));
 sky130_fd_sc_hd__and3_1 _12474_ (.A(\cur_mb_mem[162][0] ),
    .B(_06908_),
    .C(_06192_),
    .X(_07519_));
 sky130_fd_sc_hd__and3_1 _12475_ (.A(\cur_mb_mem[239][0] ),
    .B(_06149_),
    .C(_06918_),
    .X(_07520_));
 sky130_fd_sc_hd__and3_1 _12476_ (.A(\cur_mb_mem[230][0] ),
    .B(_06191_),
    .C(_06065_),
    .X(_07521_));
 sky130_fd_sc_hd__a2111o_1 _12477_ (.A1(\cur_mb_mem[56][0] ),
    .A2(_06351_),
    .B1(_07519_),
    .C1(_07520_),
    .D1(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__and3_1 _12478_ (.A(\cur_mb_mem[94][0] ),
    .B(_06895_),
    .C(_06000_),
    .X(_07523_));
 sky130_fd_sc_hd__and3_1 _12479_ (.A(\cur_mb_mem[187][0] ),
    .B(_06942_),
    .C(_06877_),
    .X(_07524_));
 sky130_fd_sc_hd__and3_1 _12480_ (.A(\cur_mb_mem[189][0] ),
    .B(_06246_),
    .C(_06216_),
    .X(_07525_));
 sky130_fd_sc_hd__a2111o_1 _12481_ (.A1(\cur_mb_mem[118][0] ),
    .A2(_06141_),
    .B1(_07523_),
    .C1(_07524_),
    .D1(_07525_),
    .X(_07526_));
 sky130_fd_sc_hd__and3_1 _12482_ (.A(\cur_mb_mem[59][0] ),
    .B(_05056_),
    .C(_06942_),
    .X(_07527_));
 sky130_fd_sc_hd__and3_1 _12483_ (.A(\cur_mb_mem[195][0] ),
    .B(_06086_),
    .C(_06091_),
    .X(_07528_));
 sky130_fd_sc_hd__and3_1 _12484_ (.A(\cur_mb_mem[99][0] ),
    .B(_06413_),
    .C(_06062_),
    .X(_07529_));
 sky130_fd_sc_hd__a2111o_1 _12485_ (.A1(\cur_mb_mem[50][0] ),
    .A2(_06172_),
    .B1(_07527_),
    .C1(_07528_),
    .D1(_07529_),
    .X(_07530_));
 sky130_fd_sc_hd__or4_2 _12486_ (.A(_07518_),
    .B(_07522_),
    .C(_07526_),
    .D(_07530_),
    .X(_07531_));
 sky130_fd_sc_hd__and3_1 _12487_ (.A(\cur_mb_mem[66][0] ),
    .B(_06380_),
    .C(_06057_),
    .X(_07532_));
 sky130_fd_sc_hd__and3_1 _12488_ (.A(\cur_mb_mem[90][0] ),
    .B(_05905_),
    .C(_07277_),
    .X(_07533_));
 sky130_fd_sc_hd__and3_1 _12489_ (.A(\cur_mb_mem[163][0] ),
    .B(_06062_),
    .C(_05922_),
    .X(_07534_));
 sky130_fd_sc_hd__a2111o_1 _12490_ (.A1(\cur_mb_mem[83][0] ),
    .A2(_06379_),
    .B1(_07532_),
    .C1(_07533_),
    .D1(_07534_),
    .X(_07535_));
 sky130_fd_sc_hd__and3_1 _12491_ (.A(\cur_mb_mem[2][0] ),
    .B(_07096_),
    .C(_06380_),
    .X(_07536_));
 sky130_fd_sc_hd__and3_1 _12492_ (.A(\cur_mb_mem[115][0] ),
    .B(_06086_),
    .C(_07253_),
    .X(_07537_));
 sky130_fd_sc_hd__and3_1 _12493_ (.A(\cur_mb_mem[147][0] ),
    .B(_06062_),
    .C(_05978_),
    .X(_07538_));
 sky130_fd_sc_hd__a2111o_1 _12494_ (.A1(\cur_mb_mem[52][0] ),
    .A2(_06241_),
    .B1(_07536_),
    .C1(_07537_),
    .D1(_07538_),
    .X(_07539_));
 sky130_fd_sc_hd__and3_1 _12495_ (.A(\cur_mb_mem[121][0] ),
    .B(_06834_),
    .C(_07253_),
    .X(_07540_));
 sky130_fd_sc_hd__and3_1 _12496_ (.A(\cur_mb_mem[140][0] ),
    .B(_06920_),
    .C(_05935_),
    .X(_07541_));
 sky130_fd_sc_hd__and3_1 _12497_ (.A(\cur_mb_mem[178][0] ),
    .B(_07099_),
    .C(_06036_),
    .X(_07542_));
 sky130_fd_sc_hd__a2111o_1 _12498_ (.A1(\cur_mb_mem[104][0] ),
    .A2(_05985_),
    .B1(_07540_),
    .C1(_07541_),
    .D1(_07542_),
    .X(_07543_));
 sky130_fd_sc_hd__and3_1 _12499_ (.A(\cur_mb_mem[18][0] ),
    .B(_07099_),
    .C(_06001_),
    .X(_07544_));
 sky130_fd_sc_hd__and3_1 _12500_ (.A(\cur_mb_mem[5][0] ),
    .B(_06112_),
    .C(_07279_),
    .X(_07545_));
 sky130_fd_sc_hd__and3_1 _12501_ (.A(\cur_mb_mem[153][0] ),
    .B(_05893_),
    .C(_05978_),
    .X(_07546_));
 sky130_fd_sc_hd__a2111o_1 _12502_ (.A1(\cur_mb_mem[30][0] ),
    .A2(_06002_),
    .B1(_07544_),
    .C1(_07545_),
    .D1(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__or4_4 _12503_ (.A(_07535_),
    .B(_07539_),
    .C(_07543_),
    .D(_07547_),
    .X(_07548_));
 sky130_fd_sc_hd__or4_1 _12504_ (.A(_07497_),
    .B(_07514_),
    .C(_07531_),
    .D(_07548_),
    .X(_07549_));
 sky130_fd_sc_hd__or4_4 _12505_ (.A(_07373_),
    .B(_07408_),
    .C(_07479_),
    .D(_07549_),
    .X(_07550_));
 sky130_fd_sc_hd__o22ai_4 _12506_ (.A1(\cur_mb_mem[0][0] ),
    .A2(_05908_),
    .B1(_07303_),
    .B2(_07550_),
    .Y(_07551_));
 sky130_fd_sc_hd__a22o_1 _12507_ (.A1(net98),
    .A2(_07286_),
    .B1(_07551_),
    .B2(net97),
    .X(_07552_));
 sky130_fd_sc_hd__or2_1 _12508_ (.A(net98),
    .B(_07286_),
    .X(_07553_));
 sky130_fd_sc_hd__a22o_1 _12509_ (.A1(\cur_mb_mem[223][3] ),
    .A2(_06151_),
    .B1(_06297_),
    .B2(\cur_mb_mem[95][3] ),
    .X(_07554_));
 sky130_fd_sc_hd__a22o_1 _12510_ (.A1(\cur_mb_mem[38][3] ),
    .A2(_06396_),
    .B1(_06075_),
    .B2(\cur_mb_mem[128][3] ),
    .X(_07555_));
 sky130_fd_sc_hd__and3_1 _12511_ (.A(\cur_mb_mem[214][3] ),
    .B(_06186_),
    .C(_05948_),
    .X(_07556_));
 sky130_fd_sc_hd__a31o_4 _12512_ (.A1(\cur_mb_mem[221][3] ),
    .A2(_05946_),
    .A3(_05942_),
    .B1(_07556_),
    .X(_07557_));
 sky130_fd_sc_hd__a211o_1 _12513_ (.A1(\cur_mb_mem[159][3] ),
    .A2(_06174_),
    .B1(_07555_),
    .C1(_07557_),
    .X(_07558_));
 sky130_fd_sc_hd__a221o_1 _12514_ (.A1(\cur_mb_mem[101][3] ),
    .A2(_06269_),
    .B1(_06242_),
    .B2(\cur_mb_mem[22][3] ),
    .C1(_07558_),
    .X(_07559_));
 sky130_fd_sc_hd__a32o_1 _12515_ (.A1(\cur_mb_mem[160][3] ),
    .A2(_06426_),
    .A3(_05972_),
    .B1(_06489_),
    .B2(\cur_mb_mem[25][3] ),
    .X(_07560_));
 sky130_fd_sc_hd__a32o_4 _12516_ (.A1(\cur_mb_mem[148][3] ),
    .A2(_06134_),
    .A3(_05979_),
    .B1(_06322_),
    .B2(\cur_mb_mem[108][3] ),
    .X(_07561_));
 sky130_fd_sc_hd__a221o_1 _12517_ (.A1(\cur_mb_mem[12][3] ),
    .A2(_05928_),
    .B1(_06193_),
    .B2(\cur_mb_mem[166][3] ),
    .C1(_07561_),
    .X(_07562_));
 sky130_fd_sc_hd__a32o_1 _12518_ (.A1(\cur_mb_mem[20][3] ),
    .A2(_06223_),
    .A3(_05976_),
    .B1(_06017_),
    .B2(\cur_mb_mem[28][3] ),
    .X(_07563_));
 sky130_fd_sc_hd__a32o_4 _12519_ (.A1(\cur_mb_mem[219][3] ),
    .A2(_06261_),
    .A3(_05948_),
    .B1(_06040_),
    .B2(\cur_mb_mem[185][3] ),
    .X(_07564_));
 sky130_fd_sc_hd__a22o_1 _12520_ (.A1(\cur_mb_mem[46][3] ),
    .A2(_06107_),
    .B1(_05966_),
    .B2(\cur_mb_mem[129][3] ),
    .X(_07565_));
 sky130_fd_sc_hd__a22o_1 _12521_ (.A1(\cur_mb_mem[45][3] ),
    .A2(_06491_),
    .B1(_06316_),
    .B2(\cur_mb_mem[176][3] ),
    .X(_07566_));
 sky130_fd_sc_hd__a32o_1 _12522_ (.A1(\cur_mb_mem[201][3] ),
    .A2(_05910_),
    .A3(_06092_),
    .B1(_06217_),
    .B2(\cur_mb_mem[180][3] ),
    .X(_07567_));
 sky130_fd_sc_hd__or4_1 _12523_ (.A(_07564_),
    .B(_07565_),
    .C(_07566_),
    .D(_07567_),
    .X(_07568_));
 sky130_fd_sc_hd__or4_1 _12524_ (.A(_07560_),
    .B(_07562_),
    .C(_07563_),
    .D(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__a2111o_2 _12525_ (.A1(\cur_mb_mem[31][3] ),
    .A2(_06178_),
    .B1(_07554_),
    .C1(_07559_),
    .D1(_07569_),
    .X(_07570_));
 sky130_fd_sc_hd__and3_1 _12526_ (.A(\cur_mb_mem[170][3] ),
    .B(_06442_),
    .C(_06333_),
    .X(_07571_));
 sky130_fd_sc_hd__and3_1 _12527_ (.A(\cur_mb_mem[81][3] ),
    .B(_06008_),
    .C(_06076_),
    .X(_07572_));
 sky130_fd_sc_hd__and3_1 _12528_ (.A(\cur_mb_mem[105][3] ),
    .B(_06038_),
    .C(_06313_),
    .X(_07573_));
 sky130_fd_sc_hd__a2111o_2 _12529_ (.A1(\cur_mb_mem[36][3] ),
    .A2(_06360_),
    .B1(_07571_),
    .C1(_07572_),
    .D1(_07573_),
    .X(_07574_));
 sky130_fd_sc_hd__and3_1 _12530_ (.A(\cur_mb_mem[89][3] ),
    .B(_05909_),
    .C(_06008_),
    .X(_07575_));
 sky130_fd_sc_hd__and3_2 _12531_ (.A(\cur_mb_mem[27][3] ),
    .B(_06003_),
    .C(_06403_),
    .X(_07576_));
 sky130_fd_sc_hd__and3_1 _12532_ (.A(\cur_mb_mem[194][3] ),
    .B(_06341_),
    .C(_06456_),
    .X(_07577_));
 sky130_fd_sc_hd__a2111o_1 _12533_ (.A1(\cur_mb_mem[141][3] ),
    .A2(_06250_),
    .B1(_07575_),
    .C1(_07576_),
    .D1(_07577_),
    .X(_07578_));
 sky130_fd_sc_hd__and3_1 _12534_ (.A(\cur_mb_mem[122][3] ),
    .B(_06442_),
    .C(_06731_),
    .X(_07579_));
 sky130_fd_sc_hd__and3_1 _12535_ (.A(\cur_mb_mem[125][3] ),
    .B(_06011_),
    .C(_06731_),
    .X(_07580_));
 sky130_fd_sc_hd__and3_1 _12536_ (.A(\cur_mb_mem[222][3] ),
    .B(_06270_),
    .C(_06435_),
    .X(_07581_));
 sky130_fd_sc_hd__a2111o_4 _12537_ (.A1(\cur_mb_mem[10][3] ),
    .A2(_06408_),
    .B1(_07579_),
    .C1(_07580_),
    .D1(_07581_),
    .X(_07582_));
 sky130_fd_sc_hd__and3_1 _12538_ (.A(\cur_mb_mem[217][3] ),
    .B(_06038_),
    .C(_06348_),
    .X(_07583_));
 sky130_fd_sc_hd__and3_1 _12539_ (.A(\cur_mb_mem[154][3] ),
    .B(_06115_),
    .C(_06434_),
    .X(_07584_));
 sky130_fd_sc_hd__and3_1 _12540_ (.A(\cur_mb_mem[124][3] ),
    .B(_06754_),
    .C(_06207_),
    .X(_07585_));
 sky130_fd_sc_hd__a2111o_2 _12541_ (.A1(\cur_mb_mem[190][3] ),
    .A2(_06480_),
    .B1(_07583_),
    .C1(_07584_),
    .D1(_07585_),
    .X(_07586_));
 sky130_fd_sc_hd__or4_1 _12542_ (.A(_07574_),
    .B(_07578_),
    .C(_07582_),
    .D(_07586_),
    .X(_07587_));
 sky130_fd_sc_hd__and3_1 _12543_ (.A(\cur_mb_mem[57][3] ),
    .B(_06849_),
    .C(_05909_),
    .X(_07588_));
 sky130_fd_sc_hd__and3_1 _12544_ (.A(\cur_mb_mem[86][3] ),
    .B(_06008_),
    .C(_06159_),
    .X(_07589_));
 sky130_fd_sc_hd__and3_1 _12545_ (.A(\cur_mb_mem[136][3] ),
    .B(_05895_),
    .C(_06382_),
    .X(_07590_));
 sky130_fd_sc_hd__a2111o_1 _12546_ (.A1(\cur_mb_mem[4][3] ),
    .A2(_06162_),
    .B1(_07588_),
    .C1(_07589_),
    .D1(_07590_),
    .X(_07591_));
 sky130_fd_sc_hd__and3_4 _12547_ (.A(\cur_mb_mem[192][3] ),
    .B(_06986_),
    .C(_06074_),
    .X(_07592_));
 sky130_fd_sc_hd__and3_1 _12548_ (.A(\cur_mb_mem[77][3] ),
    .B(_06011_),
    .C(_06428_),
    .X(_07593_));
 sky130_fd_sc_hd__and3_1 _12549_ (.A(\cur_mb_mem[58][3] ),
    .B(_06350_),
    .C(_05931_),
    .X(_07594_));
 sky130_fd_sc_hd__a2111o_1 _12550_ (.A1(\cur_mb_mem[132][3] ),
    .A2(net220),
    .B1(_07592_),
    .C1(_07593_),
    .D1(_07594_),
    .X(_07595_));
 sky130_fd_sc_hd__and3_1 _12551_ (.A(\cur_mb_mem[69][3] ),
    .B(_06428_),
    .C(_06131_),
    .X(_07596_));
 sky130_fd_sc_hd__and3_4 _12552_ (.A(\cur_mb_mem[51][3] ),
    .B(_06849_),
    .C(_06347_),
    .X(_07597_));
 sky130_fd_sc_hd__and3_1 _12553_ (.A(\cur_mb_mem[64][3] ),
    .B(_06233_),
    .C(_06815_),
    .X(_07598_));
 sky130_fd_sc_hd__a2111o_1 _12554_ (.A1(\cur_mb_mem[29][3] ),
    .A2(_06404_),
    .B1(_07596_),
    .C1(_07597_),
    .D1(_07598_),
    .X(_07599_));
 sky130_fd_sc_hd__and3_1 _12555_ (.A(\cur_mb_mem[70][3] ),
    .B(_06210_),
    .C(_06143_),
    .X(_07600_));
 sky130_fd_sc_hd__and3_1 _12556_ (.A(\cur_mb_mem[65][3] ),
    .B(_06121_),
    .C(_06353_),
    .X(_07601_));
 sky130_fd_sc_hd__and3_1 _12557_ (.A(\cur_mb_mem[78][3] ),
    .B(_06809_),
    .C(_07075_),
    .X(_07602_));
 sky130_fd_sc_hd__a2111o_1 _12558_ (.A1(\cur_mb_mem[19][3] ),
    .A2(_06282_),
    .B1(_07600_),
    .C1(_07601_),
    .D1(_07602_),
    .X(_07603_));
 sky130_fd_sc_hd__or4_4 _12559_ (.A(_07591_),
    .B(_07595_),
    .C(_07599_),
    .D(_07603_),
    .X(_07604_));
 sky130_fd_sc_hd__and3_1 _12560_ (.A(\cur_mb_mem[85][3] ),
    .B(_06008_),
    .C(_06131_),
    .X(_07605_));
 sky130_fd_sc_hd__and3_1 _12561_ (.A(\cur_mb_mem[171][3] ),
    .B(_06003_),
    .C(_06333_),
    .X(_07606_));
 sky130_fd_sc_hd__and3_2 _12562_ (.A(\cur_mb_mem[1][3] ),
    .B(_06300_),
    .C(_06353_),
    .X(_07607_));
 sky130_fd_sc_hd__a2111o_1 _12563_ (.A1(\cur_mb_mem[100][3] ),
    .A2(_06028_),
    .B1(_07605_),
    .C1(_07606_),
    .D1(_07607_),
    .X(_07608_));
 sky130_fd_sc_hd__and3_1 _12564_ (.A(\cur_mb_mem[116][3] ),
    .B(net260),
    .C(_06731_),
    .X(_07609_));
 sky130_fd_sc_hd__and3_1 _12565_ (.A(\cur_mb_mem[202][3] ),
    .B(_05904_),
    .C(_06789_),
    .X(_07610_));
 sky130_fd_sc_hd__and3_1 _12566_ (.A(\cur_mb_mem[252][3] ),
    .B(_04429_),
    .C(_05901_),
    .X(_07611_));
 sky130_fd_sc_hd__and3_1 _12567_ (.A(\cur_mb_mem[13][3] ),
    .B(_06365_),
    .C(_05944_),
    .X(_07612_));
 sky130_fd_sc_hd__or4_1 _12568_ (.A(_07609_),
    .B(_07610_),
    .C(_07611_),
    .D(_07612_),
    .X(_07613_));
 sky130_fd_sc_hd__and3_1 _12569_ (.A(\cur_mb_mem[181][3] ),
    .B(_06013_),
    .C(_06131_),
    .X(_07614_));
 sky130_fd_sc_hd__and3_1 _12570_ (.A(\cur_mb_mem[209][3] ),
    .B(_06348_),
    .C(_05995_),
    .X(_07615_));
 sky130_fd_sc_hd__and3_1 _12571_ (.A(\cur_mb_mem[200][3] ),
    .B(_06455_),
    .C(_06352_),
    .X(_07616_));
 sky130_fd_sc_hd__a2111o_2 _12572_ (.A1(\cur_mb_mem[14][3] ),
    .A2(_06367_),
    .B1(_07614_),
    .C1(_07615_),
    .D1(_07616_),
    .X(_07617_));
 sky130_fd_sc_hd__and3_1 _12573_ (.A(\cur_mb_mem[165][3] ),
    .B(_06758_),
    .C(_06220_),
    .X(_07618_));
 sky130_fd_sc_hd__and3_1 _12574_ (.A(\cur_mb_mem[126][3] ),
    .B(_06138_),
    .C(_07075_),
    .X(_07619_));
 sky130_fd_sc_hd__and3_1 _12575_ (.A(\cur_mb_mem[73][3] ),
    .B(_06903_),
    .C(_06057_),
    .X(_07620_));
 sky130_fd_sc_hd__a2111o_2 _12576_ (.A1(\cur_mb_mem[67][3] ),
    .A2(_06429_),
    .B1(_07618_),
    .C1(_07619_),
    .D1(_07620_),
    .X(_07621_));
 sky130_fd_sc_hd__or4_1 _12577_ (.A(_07608_),
    .B(_07613_),
    .C(_07617_),
    .D(_07621_),
    .X(_07622_));
 sky130_fd_sc_hd__and3_1 _12578_ (.A(\cur_mb_mem[9][3] ),
    .B(_06365_),
    .C(_06038_),
    .X(_07623_));
 sky130_fd_sc_hd__and3_1 _12579_ (.A(\cur_mb_mem[145][3] ),
    .B(_06434_),
    .C(_06353_),
    .X(_07624_));
 sky130_fd_sc_hd__and3_1 _12580_ (.A(\cur_mb_mem[158][3] ),
    .B(_06747_),
    .C(_07075_),
    .X(_07625_));
 sky130_fd_sc_hd__a2111o_2 _12581_ (.A1(\cur_mb_mem[203][3] ),
    .A2(_06325_),
    .B1(_07623_),
    .C1(_07624_),
    .D1(_07625_),
    .X(_07626_));
 sky130_fd_sc_hd__and3_1 _12582_ (.A(\cur_mb_mem[34][3] ),
    .B(_06171_),
    .C(_06395_),
    .X(_07627_));
 sky130_fd_sc_hd__and3_1 _12583_ (.A(\cur_mb_mem[186][3] ),
    .B(_06115_),
    .C(_06019_),
    .X(_07628_));
 sky130_fd_sc_hd__and3_1 _12584_ (.A(\cur_mb_mem[16][3] ),
    .B(_05970_),
    .C(_06235_),
    .X(_07629_));
 sky130_fd_sc_hd__a2111o_2 _12585_ (.A1(\cur_mb_mem[11][3] ),
    .A2(_06301_),
    .B1(_07627_),
    .C1(_07628_),
    .D1(_07629_),
    .X(_07630_));
 sky130_fd_sc_hd__and3_1 _12586_ (.A(\cur_mb_mem[35][3] ),
    .B(_06355_),
    .C(_06395_),
    .X(_07631_));
 sky130_fd_sc_hd__and3_1 _12587_ (.A(\cur_mb_mem[54][3] ),
    .B(_06856_),
    .C(_06140_),
    .X(_07632_));
 sky130_fd_sc_hd__and3_1 _12588_ (.A(\cur_mb_mem[204][3] ),
    .B(_06937_),
    .C(_06082_),
    .X(_07633_));
 sky130_fd_sc_hd__a2111o_4 _12589_ (.A1(\cur_mb_mem[131][3] ),
    .A2(_06383_),
    .B1(_07631_),
    .C1(_07632_),
    .D1(_07633_),
    .X(_07634_));
 sky130_fd_sc_hd__and3_4 _12590_ (.A(\cur_mb_mem[244][3] ),
    .B(_06165_),
    .C(_06232_),
    .X(_07635_));
 sky130_fd_sc_hd__and3_1 _12591_ (.A(\cur_mb_mem[3][3] ),
    .B(_06707_),
    .C(_06770_),
    .X(_07636_));
 sky130_fd_sc_hd__and3_1 _12592_ (.A(\cur_mb_mem[113][3] ),
    .B(_07078_),
    .C(_06251_),
    .X(_07637_));
 sky130_fd_sc_hd__a2111o_1 _12593_ (.A1(\cur_mb_mem[155][3] ),
    .A2(_06402_),
    .B1(_07635_),
    .C1(_07636_),
    .D1(_07637_),
    .X(_07638_));
 sky130_fd_sc_hd__or4_1 _12594_ (.A(_07626_),
    .B(_07630_),
    .C(_07634_),
    .D(_07638_),
    .X(_07639_));
 sky130_fd_sc_hd__or4_2 _12595_ (.A(_07587_),
    .B(_07604_),
    .C(_07622_),
    .D(_07639_),
    .X(_07640_));
 sky130_fd_sc_hd__a32o_1 _12596_ (.A1(\cur_mb_mem[247][3] ),
    .A2(_04430_),
    .A3(_06096_),
    .B1(_06248_),
    .B2(\cur_mb_mem[237][3] ),
    .X(_07641_));
 sky130_fd_sc_hd__a32o_1 _12597_ (.A1(\cur_mb_mem[175][3] ),
    .A2(_04423_),
    .A3(_06137_),
    .B1(_06447_),
    .B2(\cur_mb_mem[215][3] ),
    .X(_07642_));
 sky130_fd_sc_hd__a2111o_2 _12598_ (.A1(\cur_mb_mem[127][3] ),
    .A2(_06101_),
    .B1(_07641_),
    .C1(_07642_),
    .D1(_06185_),
    .X(_07643_));
 sky130_fd_sc_hd__a22o_1 _12599_ (.A1(\cur_mb_mem[242][3] ),
    .A2(_06335_),
    .B1(_06195_),
    .B2(\cur_mb_mem[164][3] ),
    .X(_07644_));
 sky130_fd_sc_hd__a221o_1 _12600_ (.A1(\cur_mb_mem[216][3] ),
    .A2(_06317_),
    .B1(_06433_),
    .B2(\cur_mb_mem[144][3] ),
    .C1(_07644_),
    .X(_07645_));
 sky130_fd_sc_hd__a22o_1 _12601_ (.A1(\cur_mb_mem[226][3] ),
    .A2(_06256_),
    .B1(_06180_),
    .B2(\cur_mb_mem[231][3] ),
    .X(_07646_));
 sky130_fd_sc_hd__a32o_1 _12602_ (.A1(\cur_mb_mem[235][3] ),
    .A2(_06261_),
    .A3(_06224_),
    .B1(_06344_),
    .B2(\cur_mb_mem[37][3] ),
    .X(_07647_));
 sky130_fd_sc_hd__and3_1 _12603_ (.A(\cur_mb_mem[15][3] ),
    .B(_06068_),
    .C(_06365_),
    .X(_07648_));
 sky130_fd_sc_hd__and3_1 _12604_ (.A(\cur_mb_mem[232][3] ),
    .B(_05895_),
    .C(_06116_),
    .X(_07649_));
 sky130_fd_sc_hd__and3_1 _12605_ (.A(\cur_mb_mem[234][3] ),
    .B(_06115_),
    .C(_06255_),
    .X(_07650_));
 sky130_fd_sc_hd__a2111o_1 _12606_ (.A1(\cur_mb_mem[134][3] ),
    .A2(_06211_),
    .B1(_07648_),
    .C1(_07649_),
    .D1(_07650_),
    .X(_07651_));
 sky130_fd_sc_hd__and3_1 _12607_ (.A(\cur_mb_mem[246][3] ),
    .B(_06158_),
    .C(_06140_),
    .X(_07652_));
 sky130_fd_sc_hd__and3_1 _12608_ (.A(\cur_mb_mem[227][3] ),
    .B(_06289_),
    .C(_06255_),
    .X(_07653_));
 sky130_fd_sc_hd__and3_2 _12609_ (.A(\cur_mb_mem[184][3] ),
    .B(_05982_),
    .C(_06830_),
    .X(_07654_));
 sky130_fd_sc_hd__a2111o_1 _12610_ (.A1(\cur_mb_mem[177][3] ),
    .A2(_06020_),
    .B1(_07652_),
    .C1(_07653_),
    .D1(_07654_),
    .X(_07655_));
 sky130_fd_sc_hd__or4_2 _12611_ (.A(_07646_),
    .B(_07647_),
    .C(_07651_),
    .D(_07655_),
    .X(_07656_));
 sky130_fd_sc_hd__and3_1 _12612_ (.A(\cur_mb_mem[172][3] ),
    .B(_06422_),
    .C(_06758_),
    .X(_07657_));
 sky130_fd_sc_hd__and3_1 _12613_ (.A(\cur_mb_mem[43][3] ),
    .B(_06312_),
    .C(_06395_),
    .X(_07658_));
 sky130_fd_sc_hd__and3_1 _12614_ (.A(\cur_mb_mem[88][3] ),
    .B(_06478_),
    .C(_06230_),
    .X(_07659_));
 sky130_fd_sc_hd__a2111o_1 _12615_ (.A1(\cur_mb_mem[61][3] ),
    .A2(_06359_),
    .B1(_07657_),
    .C1(_07658_),
    .D1(_07659_),
    .X(_07660_));
 sky130_fd_sc_hd__and3_4 _12616_ (.A(\cur_mb_mem[245][3] ),
    .B(_06158_),
    .C(_06220_),
    .X(_07661_));
 sky130_fd_sc_hd__and3_1 _12617_ (.A(\cur_mb_mem[112][3] ),
    .B(_06051_),
    .C(_06815_),
    .X(_07662_));
 sky130_fd_sc_hd__and3_2 _12618_ (.A(\cur_mb_mem[72][3] ),
    .B(_06478_),
    .C(_06809_),
    .X(_07663_));
 sky130_fd_sc_hd__a2111o_1 _12619_ (.A1(\cur_mb_mem[138][3] ),
    .A2(_05934_),
    .B1(_07661_),
    .C1(_07662_),
    .D1(_07663_),
    .X(_07664_));
 sky130_fd_sc_hd__and3_1 _12620_ (.A(\cur_mb_mem[133][3] ),
    .B(_06382_),
    .C(_06220_),
    .X(_07665_));
 sky130_fd_sc_hd__and3_1 _12621_ (.A(\cur_mb_mem[117][3] ),
    .B(_06138_),
    .C(_06147_),
    .X(_07666_));
 sky130_fd_sc_hd__and3_1 _12622_ (.A(\cur_mb_mem[120][3] ),
    .B(_05982_),
    .C(_06207_),
    .X(_07667_));
 sky130_fd_sc_hd__a2111o_1 _12623_ (.A1(\cur_mb_mem[97][3] ),
    .A2(_06077_),
    .B1(_07665_),
    .C1(_07666_),
    .D1(_07667_),
    .X(_07668_));
 sky130_fd_sc_hd__and3_1 _12624_ (.A(\cur_mb_mem[196][3] ),
    .B(_06026_),
    .C(_06789_),
    .X(_07669_));
 sky130_fd_sc_hd__and3_1 _12625_ (.A(\cur_mb_mem[198][3] ),
    .B(_06159_),
    .C(_06986_),
    .X(_07670_));
 sky130_fd_sc_hd__and3_1 _12626_ (.A(\cur_mb_mem[208][3] ),
    .B(_06802_),
    .C(_06074_),
    .X(_07671_));
 sky130_fd_sc_hd__and3_4 _12627_ (.A(\cur_mb_mem[75][3] ),
    .B(_06003_),
    .C(_06428_),
    .X(_07672_));
 sky130_fd_sc_hd__or4_4 _12628_ (.A(_07669_),
    .B(_07670_),
    .C(_07671_),
    .D(_07672_),
    .X(_07673_));
 sky130_fd_sc_hd__or4_4 _12629_ (.A(_07660_),
    .B(_07664_),
    .C(_07668_),
    .D(_07673_),
    .X(_07674_));
 sky130_fd_sc_hd__or4_2 _12630_ (.A(_07643_),
    .B(_07645_),
    .C(_07656_),
    .D(_07674_),
    .X(_07675_));
 sky130_fd_sc_hd__and3_1 _12631_ (.A(\cur_mb_mem[169][3] ),
    .B(_05909_),
    .C(_06333_),
    .X(_07676_));
 sky130_fd_sc_hd__and3_1 _12632_ (.A(\cur_mb_mem[168][3] ),
    .B(_05895_),
    .C(_06333_),
    .X(_07677_));
 sky130_fd_sc_hd__and3_1 _12633_ (.A(\cur_mb_mem[33][3] ),
    .B(_06395_),
    .C(_06353_),
    .X(_07678_));
 sky130_fd_sc_hd__a2111o_1 _12634_ (.A1(\cur_mb_mem[42][3] ),
    .A2(_06441_),
    .B1(_07676_),
    .C1(_07677_),
    .D1(_07678_),
    .X(_07679_));
 sky130_fd_sc_hd__and3_1 _12635_ (.A(\cur_mb_mem[102][3] ),
    .B(_06027_),
    .C(_06159_),
    .X(_07680_));
 sky130_fd_sc_hd__and3_2 _12636_ (.A(\cur_mb_mem[193][3] ),
    .B(_06324_),
    .C(_06076_),
    .X(_07681_));
 sky130_fd_sc_hd__and3_1 _12637_ (.A(\cur_mb_mem[96][3] ),
    .B(_06045_),
    .C(_06815_),
    .X(_07682_));
 sky130_fd_sc_hd__a2111o_1 _12638_ (.A1(\cur_mb_mem[74][3] ),
    .A2(_06417_),
    .B1(_07680_),
    .C1(_07681_),
    .D1(_07682_),
    .X(_07683_));
 sky130_fd_sc_hd__and3_2 _12639_ (.A(\cur_mb_mem[218][3] ),
    .B(_05931_),
    .C(_06802_),
    .X(_07684_));
 sky130_fd_sc_hd__and3_1 _12640_ (.A(\cur_mb_mem[137][3] ),
    .B(_06038_),
    .C(_06382_),
    .X(_07685_));
 sky130_fd_sc_hd__and3_1 _12641_ (.A(\cur_mb_mem[179][3] ),
    .B(_06289_),
    .C(_06760_),
    .X(_07686_));
 sky130_fd_sc_hd__a2111o_1 _12642_ (.A1(\cur_mb_mem[152][3] ),
    .A2(_06394_),
    .B1(_07684_),
    .C1(_07685_),
    .D1(_07686_),
    .X(_07687_));
 sky130_fd_sc_hd__and3_1 _12643_ (.A(\cur_mb_mem[109][3] ),
    .B(_06313_),
    .C(_06011_),
    .X(_07688_));
 sky130_fd_sc_hd__and3_1 _12644_ (.A(\cur_mb_mem[84][3] ),
    .B(_06166_),
    .C(_06931_),
    .X(_07689_));
 sky130_fd_sc_hd__and3_1 _12645_ (.A(\cur_mb_mem[251][3] ),
    .B(_06916_),
    .C(_06387_),
    .X(_07690_));
 sky130_fd_sc_hd__a2111o_1 _12646_ (.A1(\cur_mb_mem[110][3] ),
    .A2(_06047_),
    .B1(_07688_),
    .C1(_07689_),
    .D1(_07690_),
    .X(_07691_));
 sky130_fd_sc_hd__or4_4 _12647_ (.A(_07679_),
    .B(_07683_),
    .C(_07687_),
    .D(_07691_),
    .X(_07692_));
 sky130_fd_sc_hd__and3_1 _12648_ (.A(\cur_mb_mem[80][3] ),
    .B(_06008_),
    .C(_06074_),
    .X(_07693_));
 sky130_fd_sc_hd__and3_1 _12649_ (.A(\cur_mb_mem[17][3] ),
    .B(_06076_),
    .C(_06488_),
    .X(_07694_));
 sky130_fd_sc_hd__and3_1 _12650_ (.A(\cur_mb_mem[62][3] ),
    .B(_06350_),
    .C(_06435_),
    .X(_07695_));
 sky130_fd_sc_hd__a2111o_2 _12651_ (.A1(\cur_mb_mem[24][3] ),
    .A2(_06285_),
    .B1(_07693_),
    .C1(_07694_),
    .D1(_07695_),
    .X(_07696_));
 sky130_fd_sc_hd__and3_1 _12652_ (.A(\cur_mb_mem[130][3] ),
    .B(_06079_),
    .C(_05933_),
    .X(_07697_));
 sky130_fd_sc_hd__and3_4 _12653_ (.A(\cur_mb_mem[197][3] ),
    .B(_06324_),
    .C(_06131_),
    .X(_07698_));
 sky130_fd_sc_hd__and3_1 _12654_ (.A(\cur_mb_mem[92][3] ),
    .B(_06718_),
    .C(_06378_),
    .X(_07699_));
 sky130_fd_sc_hd__a2111o_1 _12655_ (.A1(\cur_mb_mem[161][3] ),
    .A2(_06334_),
    .B1(_07697_),
    .C1(_07698_),
    .D1(_07699_),
    .X(_07700_));
 sky130_fd_sc_hd__and3_1 _12656_ (.A(\cur_mb_mem[106][3] ),
    .B(_05931_),
    .C(_06313_),
    .X(_07701_));
 sky130_fd_sc_hd__and3_1 _12657_ (.A(\cur_mb_mem[188][3] ),
    .B(_06422_),
    .C(_06039_),
    .X(_07702_));
 sky130_fd_sc_hd__and3_1 _12658_ (.A(\cur_mb_mem[82][3] ),
    .B(_06254_),
    .C(_05914_),
    .X(_07703_));
 sky130_fd_sc_hd__a2111o_1 _12659_ (.A1(\cur_mb_mem[44][3] ),
    .A2(_06399_),
    .B1(_07701_),
    .C1(_07702_),
    .D1(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__and3_1 _12660_ (.A(\cur_mb_mem[254][3] ),
    .B(_06158_),
    .C(_06435_),
    .X(_07705_));
 sky130_fd_sc_hd__and3_1 _12661_ (.A(\cur_mb_mem[150][3] ),
    .B(_06204_),
    .C(_06434_),
    .X(_07706_));
 sky130_fd_sc_hd__and3_1 _12662_ (.A(\cur_mb_mem[212][3] ),
    .B(_06215_),
    .C(_06150_),
    .X(_07707_));
 sky130_fd_sc_hd__a2111o_4 _12663_ (.A1(\cur_mb_mem[253][3] ),
    .A2(_06034_),
    .B1(_07705_),
    .C1(_07706_),
    .D1(_07707_),
    .X(_07708_));
 sky130_fd_sc_hd__or4_2 _12664_ (.A(_07696_),
    .B(_07700_),
    .C(_07704_),
    .D(_07708_),
    .X(_07709_));
 sky130_fd_sc_hd__and3_1 _12665_ (.A(\cur_mb_mem[93][3] ),
    .B(_05913_),
    .C(_05944_),
    .X(_07710_));
 sky130_fd_sc_hd__and3_1 _12666_ (.A(\cur_mb_mem[220][3] ),
    .B(_05901_),
    .C(_05940_),
    .X(_07711_));
 sky130_fd_sc_hd__and3_1 _12667_ (.A(\cur_mb_mem[174][3] ),
    .B(_05953_),
    .C(_05921_),
    .X(_07712_));
 sky130_fd_sc_hd__and3_1 _12668_ (.A(\cur_mb_mem[206][3] ),
    .B(_05953_),
    .C(_06789_),
    .X(_07713_));
 sky130_fd_sc_hd__or4_1 _12669_ (.A(_07710_),
    .B(_07711_),
    .C(_07712_),
    .D(_07713_),
    .X(_07714_));
 sky130_fd_sc_hd__and3_2 _12670_ (.A(\cur_mb_mem[32][3] ),
    .B(_06005_),
    .C(_06009_),
    .X(_07715_));
 sky130_fd_sc_hd__and3_1 _12671_ (.A(\cur_mb_mem[8][3] ),
    .B(_06365_),
    .C(_05895_),
    .X(_07716_));
 sky130_fd_sc_hd__and3_1 _12672_ (.A(\cur_mb_mem[156][3] ),
    .B(_06754_),
    .C(_06401_),
    .X(_07717_));
 sky130_fd_sc_hd__a2111o_1 _12673_ (.A1(\cur_mb_mem[211][3] ),
    .A2(_06349_),
    .B1(_07715_),
    .C1(_07716_),
    .D1(_07717_),
    .X(_07718_));
 sky130_fd_sc_hd__and3_1 _12674_ (.A(\cur_mb_mem[157][3] ),
    .B(_06011_),
    .C(_06434_),
    .X(_07719_));
 sky130_fd_sc_hd__and3_1 _12675_ (.A(\cur_mb_mem[21][3] ),
    .B(_06475_),
    .C(_06220_),
    .X(_07720_));
 sky130_fd_sc_hd__and3_1 _12676_ (.A(\cur_mb_mem[249][3] ),
    .B(_06165_),
    .C(_06723_),
    .X(_07721_));
 sky130_fd_sc_hd__a2111o_1 _12677_ (.A1(\cur_mb_mem[250][3] ),
    .A2(_06443_),
    .B1(_07719_),
    .C1(_07720_),
    .D1(_07721_),
    .X(_07722_));
 sky130_fd_sc_hd__and3_1 _12678_ (.A(\cur_mb_mem[213][3] ),
    .B(_06270_),
    .C(_06812_),
    .X(_07723_));
 sky130_fd_sc_hd__and3_1 _12679_ (.A(\cur_mb_mem[149][3] ),
    .B(_06401_),
    .C(_06147_),
    .X(_07724_));
 sky130_fd_sc_hd__and3_1 _12680_ (.A(\cur_mb_mem[107][3] ),
    .B(_06387_),
    .C(_06268_),
    .X(_07725_));
 sky130_fd_sc_hd__a2111o_1 _12681_ (.A1(\cur_mb_mem[6][3] ),
    .A2(_06203_),
    .B1(_07723_),
    .C1(_07724_),
    .D1(_07725_),
    .X(_07726_));
 sky130_fd_sc_hd__or4_4 _12682_ (.A(_07714_),
    .B(_07718_),
    .C(_07722_),
    .D(_07726_),
    .X(_07727_));
 sky130_fd_sc_hd__and3_1 _12683_ (.A(\cur_mb_mem[243][3] ),
    .B(_06158_),
    .C(_06355_),
    .X(_07728_));
 sky130_fd_sc_hd__and3_1 _12684_ (.A(\cur_mb_mem[229][3] ),
    .B(_06812_),
    .C(_06255_),
    .X(_07729_));
 sky130_fd_sc_hd__and3_1 _12685_ (.A(\cur_mb_mem[60][3] ),
    .B(_06198_),
    .C(_06937_),
    .X(_07730_));
 sky130_fd_sc_hd__a2111o_2 _12686_ (.A1(\cur_mb_mem[53][3] ),
    .A2(_06221_),
    .B1(_07728_),
    .C1(_07729_),
    .D1(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__and3_1 _12687_ (.A(\cur_mb_mem[207][3] ),
    .B(_06120_),
    .C(_06456_),
    .X(_07732_));
 sky130_fd_sc_hd__and3_1 _12688_ (.A(\cur_mb_mem[236][3] ),
    .B(_06718_),
    .C(_06255_),
    .X(_07733_));
 sky130_fd_sc_hd__and3_1 _12689_ (.A(\cur_mb_mem[167][3] ),
    .B(_06192_),
    .C(_06708_),
    .X(_07734_));
 sky130_fd_sc_hd__a2111o_1 _12690_ (.A1(\cur_mb_mem[79][3] ),
    .A2(_06122_),
    .B1(_07732_),
    .C1(_07733_),
    .D1(_07734_),
    .X(_07735_));
 sky130_fd_sc_hd__and3_1 _12691_ (.A(\cur_mb_mem[48][3] ),
    .B(_06856_),
    .C(_06815_),
    .X(_07736_));
 sky130_fd_sc_hd__and3_1 _12692_ (.A(\cur_mb_mem[241][3] ),
    .B(_06165_),
    .C(_06841_),
    .X(_07737_));
 sky130_fd_sc_hd__and3_1 _12693_ (.A(\cur_mb_mem[41][3] ),
    .B(_06834_),
    .C(_06087_),
    .X(_07738_));
 sky130_fd_sc_hd__a2111o_1 _12694_ (.A1(\cur_mb_mem[182][3] ),
    .A2(_06205_),
    .B1(_07736_),
    .C1(_07737_),
    .D1(_07738_),
    .X(_07739_));
 sky130_fd_sc_hd__and3_1 _12695_ (.A(\cur_mb_mem[26][3] ),
    .B(_06442_),
    .C(net2006),
    .X(_07740_));
 sky130_fd_sc_hd__and3_1 _12696_ (.A(\cur_mb_mem[240][3] ),
    .B(_06032_),
    .C(_06074_),
    .X(_07741_));
 sky130_fd_sc_hd__and3_1 _12697_ (.A(\cur_mb_mem[183][3] ),
    .B(_06013_),
    .C(_06851_),
    .X(_07742_));
 sky130_fd_sc_hd__and3_2 _12698_ (.A(\cur_mb_mem[23][3] ),
    .B(_06461_),
    .C(_06488_),
    .X(_07743_));
 sky130_fd_sc_hd__or4_1 _12699_ (.A(_07740_),
    .B(_07741_),
    .C(_07742_),
    .D(_07743_),
    .X(_07744_));
 sky130_fd_sc_hd__or4_4 _12700_ (.A(_07731_),
    .B(_07735_),
    .C(_07739_),
    .D(_07744_),
    .X(_07745_));
 sky130_fd_sc_hd__or4_2 _12701_ (.A(_07692_),
    .B(_07709_),
    .C(_07727_),
    .D(_07745_),
    .X(_07746_));
 sky130_fd_sc_hd__and3_1 _12702_ (.A(\cur_mb_mem[63][3] ),
    .B(_06068_),
    .C(_06170_),
    .X(_07747_));
 sky130_fd_sc_hd__and3_1 _12703_ (.A(\cur_mb_mem[224][3] ),
    .B(_06009_),
    .C(_06116_),
    .X(_07748_));
 sky130_fd_sc_hd__and3_1 _12704_ (.A(\cur_mb_mem[191][3] ),
    .B(_06466_),
    .C(_06760_),
    .X(_07749_));
 sky130_fd_sc_hd__a2111o_4 _12705_ (.A1(\cur_mb_mem[255][3] ),
    .A2(_06304_),
    .B1(_07747_),
    .C1(_07748_),
    .D1(_07749_),
    .X(_07750_));
 sky130_fd_sc_hd__and3_1 _12706_ (.A(\cur_mb_mem[111][3] ),
    .B(_06099_),
    .C(_06267_),
    .X(_07751_));
 sky130_fd_sc_hd__and3_1 _12707_ (.A(\cur_mb_mem[71][3] ),
    .B(_06022_),
    .C(_06851_),
    .X(_07752_));
 sky130_fd_sc_hd__and3_1 _12708_ (.A(\cur_mb_mem[103][3] ),
    .B(_06267_),
    .C(_06851_),
    .X(_07753_));
 sky130_fd_sc_hd__and3_1 _12709_ (.A(\cur_mb_mem[47][3] ),
    .B(_06099_),
    .C(_06005_),
    .X(_07754_));
 sky130_fd_sc_hd__or4_4 _12710_ (.A(_07751_),
    .B(_07752_),
    .C(_07753_),
    .D(_07754_),
    .X(_07755_));
 sky130_fd_sc_hd__and3_1 _12711_ (.A(\cur_mb_mem[40][3] ),
    .B(_06455_),
    .C(_06395_),
    .X(_07756_));
 sky130_fd_sc_hd__and3_1 _12712_ (.A(\cur_mb_mem[98][3] ),
    .B(_06341_),
    .C(_05984_),
    .X(_07757_));
 sky130_fd_sc_hd__and3_1 _12713_ (.A(\cur_mb_mem[210][3] ),
    .B(_06080_),
    .C(_06150_),
    .X(_07758_));
 sky130_fd_sc_hd__a2111o_1 _12714_ (.A1(\cur_mb_mem[91][3] ),
    .A2(_06361_),
    .B1(_07756_),
    .C1(_07757_),
    .D1(_07758_),
    .X(_07759_));
 sky130_fd_sc_hd__and3_4 _12715_ (.A(\cur_mb_mem[238][3] ),
    .B(_07075_),
    .C(_06766_),
    .X(_07760_));
 sky130_fd_sc_hd__and3_1 _12716_ (.A(\cur_mb_mem[151][3] ),
    .B(_06747_),
    .C(_06708_),
    .X(_07761_));
 sky130_fd_sc_hd__and3_1 _12717_ (.A(\cur_mb_mem[123][3] ),
    .B(_06942_),
    .C(_07078_),
    .X(_07762_));
 sky130_fd_sc_hd__a2111o_1 _12718_ (.A1(\cur_mb_mem[68][3] ),
    .A2(_06234_),
    .B1(_07760_),
    .C1(_07761_),
    .D1(_07762_),
    .X(_07763_));
 sky130_fd_sc_hd__or4_4 _12719_ (.A(_07750_),
    .B(_07755_),
    .C(_07759_),
    .D(_07763_),
    .X(_07764_));
 sky130_fd_sc_hd__and3_4 _12720_ (.A(\cur_mb_mem[146][3] ),
    .B(_06171_),
    .C(_06434_),
    .X(_07765_));
 sky130_fd_sc_hd__and3_1 _12721_ (.A(\cur_mb_mem[199][3] ),
    .B(_06456_),
    .C(_06179_),
    .X(_07766_));
 sky130_fd_sc_hd__and3_1 _12722_ (.A(\cur_mb_mem[87][3] ),
    .B(_06230_),
    .C(_06372_),
    .X(_07767_));
 sky130_fd_sc_hd__a2111o_1 _12723_ (.A1(\cur_mb_mem[135][3] ),
    .A2(_06462_),
    .B1(_07765_),
    .C1(_07766_),
    .D1(_07767_),
    .X(_07768_));
 sky130_fd_sc_hd__and3_2 _12724_ (.A(\cur_mb_mem[76][3] ),
    .B(_06422_),
    .C(_06121_),
    .X(_07769_));
 sky130_fd_sc_hd__and3_4 _12725_ (.A(\cur_mb_mem[114][3] ),
    .B(_06341_),
    .C(_06051_),
    .X(_07770_));
 sky130_fd_sc_hd__and3_1 _12726_ (.A(\cur_mb_mem[49][3] ),
    .B(_06240_),
    .C(_06912_),
    .X(_07771_));
 sky130_fd_sc_hd__a2111o_1 _12727_ (.A1(\cur_mb_mem[225][3] ),
    .A2(_05998_),
    .B1(_07769_),
    .C1(_07770_),
    .D1(_07771_),
    .X(_07772_));
 sky130_fd_sc_hd__and3_1 _12728_ (.A(\cur_mb_mem[7][3] ),
    .B(_06300_),
    .C(_06179_),
    .X(_07773_));
 sky130_fd_sc_hd__and3_4 _12729_ (.A(\cur_mb_mem[119][3] ),
    .B(_06138_),
    .C(_06372_),
    .X(_07774_));
 sky130_fd_sc_hd__and3_1 _12730_ (.A(\cur_mb_mem[233][3] ),
    .B(_06903_),
    .C(_06247_),
    .X(_07775_));
 sky130_fd_sc_hd__a2111o_1 _12731_ (.A1(\cur_mb_mem[248][3] ),
    .A2(_06411_),
    .B1(_07773_),
    .C1(_07774_),
    .D1(_07775_),
    .X(_07776_));
 sky130_fd_sc_hd__and3_1 _12732_ (.A(\cur_mb_mem[55][3] ),
    .B(_06856_),
    .C(_06372_),
    .X(_07777_));
 sky130_fd_sc_hd__and3_1 _12733_ (.A(\cur_mb_mem[143][3] ),
    .B(_06149_),
    .C(_06146_),
    .X(_07778_));
 sky130_fd_sc_hd__and3_1 _12734_ (.A(\cur_mb_mem[228][3] ),
    .B(_06215_),
    .C(_06918_),
    .X(_07779_));
 sky130_fd_sc_hd__a2111o_1 _12735_ (.A1(\cur_mb_mem[39][3] ),
    .A2(_06373_),
    .B1(_07777_),
    .C1(_07778_),
    .D1(_07779_),
    .X(_07780_));
 sky130_fd_sc_hd__or4_2 _12736_ (.A(_07768_),
    .B(_07772_),
    .C(_07776_),
    .D(_07780_),
    .X(_07781_));
 sky130_fd_sc_hd__and3_1 _12737_ (.A(\cur_mb_mem[173][3] ),
    .B(_06011_),
    .C(_06758_),
    .X(_07782_));
 sky130_fd_sc_hd__and3_1 _12738_ (.A(\cur_mb_mem[205][3] ),
    .B(_06490_),
    .C(_06352_),
    .X(_07783_));
 sky130_fd_sc_hd__and3_1 _12739_ (.A(\cur_mb_mem[139][3] ),
    .B(_06400_),
    .C(_06146_),
    .X(_07784_));
 sky130_fd_sc_hd__a2111o_2 _12740_ (.A1(\cur_mb_mem[142][3] ),
    .A2(_06487_),
    .B1(_07782_),
    .C1(_07783_),
    .D1(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__and3_1 _12741_ (.A(\cur_mb_mem[162][3] ),
    .B(_06341_),
    .C(_06758_),
    .X(_07786_));
 sky130_fd_sc_hd__and3_1 _12742_ (.A(\cur_mb_mem[239][3] ),
    .B(_06466_),
    .C(_06255_),
    .X(_07787_));
 sky130_fd_sc_hd__and3_1 _12743_ (.A(\cur_mb_mem[230][3] ),
    .B(_06199_),
    .C(_06247_),
    .X(_07788_));
 sky130_fd_sc_hd__a2111o_1 _12744_ (.A1(\cur_mb_mem[56][3] ),
    .A2(_06351_),
    .B1(_07786_),
    .C1(_07787_),
    .D1(_07788_),
    .X(_07789_));
 sky130_fd_sc_hd__and3_1 _12745_ (.A(\cur_mb_mem[94][3] ),
    .B(_06931_),
    .C(_07075_),
    .X(_07790_));
 sky130_fd_sc_hd__and3_1 _12746_ (.A(\cur_mb_mem[187][3] ),
    .B(_06474_),
    .C(_06760_),
    .X(_07791_));
 sky130_fd_sc_hd__and3_1 _12747_ (.A(\cur_mb_mem[189][3] ),
    .B(_06056_),
    .C(_06830_),
    .X(_07792_));
 sky130_fd_sc_hd__a2111o_1 _12748_ (.A1(\cur_mb_mem[118][3] ),
    .A2(_06141_),
    .B1(_07790_),
    .C1(_07791_),
    .D1(_07792_),
    .X(_07793_));
 sky130_fd_sc_hd__and3_1 _12749_ (.A(\cur_mb_mem[59][3] ),
    .B(_06240_),
    .C(_06400_),
    .X(_07794_));
 sky130_fd_sc_hd__and3_1 _12750_ (.A(\cur_mb_mem[195][3] ),
    .B(_06980_),
    .C(_06967_),
    .X(_07795_));
 sky130_fd_sc_hd__and3_1 _12751_ (.A(\cur_mb_mem[99][3] ),
    .B(_06413_),
    .C(_06086_),
    .X(_07796_));
 sky130_fd_sc_hd__a2111o_1 _12752_ (.A1(\cur_mb_mem[50][3] ),
    .A2(_06172_),
    .B1(_07794_),
    .C1(_07795_),
    .D1(_07796_),
    .X(_07797_));
 sky130_fd_sc_hd__or4_2 _12753_ (.A(_07785_),
    .B(_07789_),
    .C(_07793_),
    .D(_07797_),
    .X(_07798_));
 sky130_fd_sc_hd__and3_1 _12754_ (.A(\cur_mb_mem[66][3] ),
    .B(_06254_),
    .C(_06809_),
    .X(_07799_));
 sky130_fd_sc_hd__and3_1 _12755_ (.A(\cur_mb_mem[90][3] ),
    .B(_05957_),
    .C(_06927_),
    .X(_07800_));
 sky130_fd_sc_hd__and3_1 _12756_ (.A(\cur_mb_mem[163][3] ),
    .B(_06980_),
    .C(_07001_),
    .X(_07801_));
 sky130_fd_sc_hd__a2111o_1 _12757_ (.A1(\cur_mb_mem[83][3] ),
    .A2(_06379_),
    .B1(_07799_),
    .C1(_07800_),
    .D1(_07801_),
    .X(_07802_));
 sky130_fd_sc_hd__and3_1 _12758_ (.A(\cur_mb_mem[2][3] ),
    .B(_06202_),
    .C(_06254_),
    .X(_07803_));
 sky130_fd_sc_hd__and3_1 _12759_ (.A(\cur_mb_mem[115][3] ),
    .B(_06770_),
    .C(_06207_),
    .X(_07804_));
 sky130_fd_sc_hd__and3_1 _12760_ (.A(\cur_mb_mem[147][3] ),
    .B(_06980_),
    .C(_06152_),
    .X(_07805_));
 sky130_fd_sc_hd__a2111o_1 _12761_ (.A1(\cur_mb_mem[52][3] ),
    .A2(_06241_),
    .B1(_07803_),
    .C1(_07804_),
    .D1(_07805_),
    .X(_07806_));
 sky130_fd_sc_hd__and3_1 _12762_ (.A(\cur_mb_mem[121][3] ),
    .B(_06723_),
    .C(_06207_),
    .X(_07807_));
 sky130_fd_sc_hd__and3_1 _12763_ (.A(\cur_mb_mem[140][3] ),
    .B(_06937_),
    .C(_06859_),
    .X(_07808_));
 sky130_fd_sc_hd__and3_1 _12764_ (.A(\cur_mb_mem[178][3] ),
    .B(_06380_),
    .C(_06877_),
    .X(_07809_));
 sky130_fd_sc_hd__a2111o_1 _12765_ (.A1(\cur_mb_mem[104][3] ),
    .A2(_05985_),
    .B1(_07807_),
    .C1(_07808_),
    .D1(_07809_),
    .X(_07810_));
 sky130_fd_sc_hd__and3_1 _12766_ (.A(\cur_mb_mem[18][3] ),
    .B(_06908_),
    .C(_06001_),
    .X(_07811_));
 sky130_fd_sc_hd__and3_1 _12767_ (.A(\cur_mb_mem[5][3] ),
    .B(_07096_),
    .C(_07279_),
    .X(_07812_));
 sky130_fd_sc_hd__and3_2 _12768_ (.A(\cur_mb_mem[153][3] ),
    .B(_05893_),
    .C(_07100_),
    .X(_07813_));
 sky130_fd_sc_hd__a2111o_1 _12769_ (.A1(\cur_mb_mem[30][3] ),
    .A2(_06002_),
    .B1(_07811_),
    .C1(_07812_),
    .D1(_07813_),
    .X(_07814_));
 sky130_fd_sc_hd__or4_4 _12770_ (.A(_07802_),
    .B(_07806_),
    .C(_07810_),
    .D(_07814_),
    .X(_07815_));
 sky130_fd_sc_hd__or4_1 _12771_ (.A(_07764_),
    .B(_07781_),
    .C(_07798_),
    .D(_07815_),
    .X(_07816_));
 sky130_fd_sc_hd__or4_4 _12772_ (.A(_07640_),
    .B(_07675_),
    .C(_07746_),
    .D(_07816_),
    .X(_07817_));
 sky130_fd_sc_hd__o22ai_4 _12773_ (.A1(\cur_mb_mem[0][3] ),
    .A2(_05908_),
    .B1(_07570_),
    .B2(_07817_),
    .Y(_07818_));
 sky130_fd_sc_hd__xnor2_1 _12774_ (.A(net100),
    .B(_07818_),
    .Y(_07819_));
 sky130_fd_sc_hd__nor2_1 _12775_ (.A(\cur_mb_mem[0][2] ),
    .B(_05908_),
    .Y(_07820_));
 sky130_fd_sc_hd__a22o_1 _12776_ (.A1(\cur_mb_mem[223][2] ),
    .A2(_06151_),
    .B1(_06297_),
    .B2(\cur_mb_mem[95][2] ),
    .X(_07821_));
 sky130_fd_sc_hd__a22o_1 _12777_ (.A1(\cur_mb_mem[38][2] ),
    .A2(_06396_),
    .B1(_06075_),
    .B2(\cur_mb_mem[128][2] ),
    .X(_07822_));
 sky130_fd_sc_hd__and3_1 _12778_ (.A(\cur_mb_mem[214][2] ),
    .B(_06186_),
    .C(_05948_),
    .X(_07823_));
 sky130_fd_sc_hd__a31o_4 _12779_ (.A1(\cur_mb_mem[221][2] ),
    .A2(_05946_),
    .A3(_05942_),
    .B1(_07823_),
    .X(_07824_));
 sky130_fd_sc_hd__a211o_1 _12780_ (.A1(\cur_mb_mem[159][2] ),
    .A2(_06174_),
    .B1(_07822_),
    .C1(_07824_),
    .X(_07825_));
 sky130_fd_sc_hd__a221o_1 _12781_ (.A1(\cur_mb_mem[101][2] ),
    .A2(_06269_),
    .B1(_06242_),
    .B2(\cur_mb_mem[22][2] ),
    .C1(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__a32o_1 _12782_ (.A1(\cur_mb_mem[160][2] ),
    .A2(_06426_),
    .A3(_05972_),
    .B1(_06489_),
    .B2(\cur_mb_mem[25][2] ),
    .X(_07827_));
 sky130_fd_sc_hd__a32o_4 _12783_ (.A1(\cur_mb_mem[148][2] ),
    .A2(_06134_),
    .A3(_05979_),
    .B1(_06322_),
    .B2(\cur_mb_mem[108][2] ),
    .X(_07828_));
 sky130_fd_sc_hd__a221o_1 _12784_ (.A1(\cur_mb_mem[12][2] ),
    .A2(_05928_),
    .B1(_06193_),
    .B2(\cur_mb_mem[166][2] ),
    .C1(_07828_),
    .X(_07829_));
 sky130_fd_sc_hd__a32o_1 _12785_ (.A1(\cur_mb_mem[20][2] ),
    .A2(_06223_),
    .A3(_05976_),
    .B1(_06017_),
    .B2(\cur_mb_mem[28][2] ),
    .X(_07830_));
 sky130_fd_sc_hd__a32o_4 _12786_ (.A1(\cur_mb_mem[219][2] ),
    .A2(_06261_),
    .A3(_05948_),
    .B1(_06040_),
    .B2(\cur_mb_mem[185][2] ),
    .X(_07831_));
 sky130_fd_sc_hd__a22o_1 _12787_ (.A1(\cur_mb_mem[46][2] ),
    .A2(_06107_),
    .B1(_05966_),
    .B2(\cur_mb_mem[129][2] ),
    .X(_07832_));
 sky130_fd_sc_hd__a22o_1 _12788_ (.A1(\cur_mb_mem[45][2] ),
    .A2(_06491_),
    .B1(_06316_),
    .B2(\cur_mb_mem[176][2] ),
    .X(_07833_));
 sky130_fd_sc_hd__a32o_1 _12789_ (.A1(\cur_mb_mem[201][2] ),
    .A2(_05911_),
    .A3(_06092_),
    .B1(_06217_),
    .B2(\cur_mb_mem[180][2] ),
    .X(_07834_));
 sky130_fd_sc_hd__or4_1 _12790_ (.A(_07831_),
    .B(_07832_),
    .C(_07833_),
    .D(_07834_),
    .X(_07835_));
 sky130_fd_sc_hd__or4_1 _12791_ (.A(_07827_),
    .B(_07829_),
    .C(_07830_),
    .D(_07835_),
    .X(_07836_));
 sky130_fd_sc_hd__a2111o_1 _12792_ (.A1(\cur_mb_mem[31][2] ),
    .A2(_06178_),
    .B1(_07821_),
    .C1(_07826_),
    .D1(_07836_),
    .X(_07837_));
 sky130_fd_sc_hd__and3_1 _12793_ (.A(\cur_mb_mem[170][2] ),
    .B(_06035_),
    .C(_05956_),
    .X(_07838_));
 sky130_fd_sc_hd__a31o_1 _12794_ (.A1(\cur_mb_mem[105][2] ),
    .A2(_05912_),
    .A3(_06299_),
    .B1(_07838_),
    .X(_07839_));
 sky130_fd_sc_hd__a32o_1 _12795_ (.A1(\cur_mb_mem[81][2] ),
    .A2(_05916_),
    .A3(_05994_),
    .B1(_06360_),
    .B2(\cur_mb_mem[36][2] ),
    .X(_07840_));
 sky130_fd_sc_hd__a32o_1 _12796_ (.A1(\cur_mb_mem[89][2] ),
    .A2(_06336_),
    .A3(_05925_),
    .B1(_06250_),
    .B2(\cur_mb_mem[141][2] ),
    .X(_07841_));
 sky130_fd_sc_hd__a22o_1 _12797_ (.A1(\cur_mb_mem[27][2] ),
    .A2(_06476_),
    .B1(_06083_),
    .B2(\cur_mb_mem[194][2] ),
    .X(_07842_));
 sky130_fd_sc_hd__and3_1 _12798_ (.A(\cur_mb_mem[122][2] ),
    .B(_05905_),
    .C(_07021_),
    .X(_07843_));
 sky130_fd_sc_hd__and3_1 _12799_ (.A(\cur_mb_mem[125][2] ),
    .B(_05945_),
    .C(_06052_),
    .X(_07844_));
 sky130_fd_sc_hd__and3_1 _12800_ (.A(\cur_mb_mem[222][2] ),
    .B(_05941_),
    .C(_05954_),
    .X(_07845_));
 sky130_fd_sc_hd__a2111o_1 _12801_ (.A1(\cur_mb_mem[10][2] ),
    .A2(_06408_),
    .B1(_07843_),
    .C1(_07844_),
    .D1(_07845_),
    .X(_07846_));
 sky130_fd_sc_hd__and3_1 _12802_ (.A(\cur_mb_mem[154][2] ),
    .B(_05958_),
    .C(_05978_),
    .X(_07847_));
 sky130_fd_sc_hd__a31o_1 _12803_ (.A1(\cur_mb_mem[124][2] ),
    .A2(_05937_),
    .A3(_06118_),
    .B1(_07847_),
    .X(_07848_));
 sky130_fd_sc_hd__a32o_1 _12804_ (.A1(\cur_mb_mem[217][2] ),
    .A2(_05911_),
    .A3(_05948_),
    .B1(_06480_),
    .B2(\cur_mb_mem[190][2] ),
    .X(_07849_));
 sky130_fd_sc_hd__or3_4 _12805_ (.A(_07846_),
    .B(_07848_),
    .C(_07849_),
    .X(_07850_));
 sky130_fd_sc_hd__or3_2 _12806_ (.A(_07841_),
    .B(_07842_),
    .C(_07850_),
    .X(_07851_));
 sky130_fd_sc_hd__or3_2 _12807_ (.A(_07839_),
    .B(_07840_),
    .C(_07851_),
    .X(_07852_));
 sky130_fd_sc_hd__a32o_1 _12808_ (.A1(\cur_mb_mem[86][2] ),
    .A2(_05916_),
    .A3(_06187_),
    .B1(_06162_),
    .B2(\cur_mb_mem[4][2] ),
    .X(_07853_));
 sky130_fd_sc_hd__a32o_1 _12809_ (.A1(\cur_mb_mem[57][2] ),
    .A2(_05059_),
    .A3(_05912_),
    .B1(_06292_),
    .B2(\cur_mb_mem[136][2] ),
    .X(_07854_));
 sky130_fd_sc_hd__and3_1 _12810_ (.A(\cur_mb_mem[192][2] ),
    .B(_06092_),
    .C(_05971_),
    .X(_07855_));
 sky130_fd_sc_hd__a31o_1 _12811_ (.A1(\cur_mb_mem[58][2] ),
    .A2(_05058_),
    .A3(_06035_),
    .B1(_07855_),
    .X(_07856_));
 sky130_fd_sc_hd__a22o_1 _12812_ (.A1(\cur_mb_mem[132][2] ),
    .A2(net220),
    .B1(_06058_),
    .B2(\cur_mb_mem[77][2] ),
    .X(_07857_));
 sky130_fd_sc_hd__a32o_1 _12813_ (.A1(\cur_mb_mem[78][2] ),
    .A2(_06024_),
    .A3(_05954_),
    .B1(_06282_),
    .B2(\cur_mb_mem[19][2] ),
    .X(_07858_));
 sky130_fd_sc_hd__a32o_1 _12814_ (.A1(\cur_mb_mem[64][2] ),
    .A2(_06024_),
    .A3(_05971_),
    .B1(_06404_),
    .B2(\cur_mb_mem[29][2] ),
    .X(_07859_));
 sky130_fd_sc_hd__a32o_1 _12815_ (.A1(\cur_mb_mem[51][2] ),
    .A2(_05057_),
    .A3(_06063_),
    .B1(_06218_),
    .B2(\cur_mb_mem[69][2] ),
    .X(_07860_));
 sky130_fd_sc_hd__a22o_1 _12816_ (.A1(\cur_mb_mem[70][2] ),
    .A2(_06144_),
    .B1(_06483_),
    .B2(\cur_mb_mem[65][2] ),
    .X(_07861_));
 sky130_fd_sc_hd__or4_1 _12817_ (.A(_07858_),
    .B(_07859_),
    .C(_07860_),
    .D(_07861_),
    .X(_07862_));
 sky130_fd_sc_hd__or3_1 _12818_ (.A(_07856_),
    .B(_07857_),
    .C(_07862_),
    .X(_07863_));
 sky130_fd_sc_hd__a32o_2 _12819_ (.A1(\cur_mb_mem[16][2] ),
    .A2(_05971_),
    .A3(_05975_),
    .B1(_06301_),
    .B2(\cur_mb_mem[11][2] ),
    .X(_07864_));
 sky130_fd_sc_hd__a22o_1 _12820_ (.A1(\cur_mb_mem[203][2] ),
    .A2(_06325_),
    .B1(_06252_),
    .B2(\cur_mb_mem[145][2] ),
    .X(_07865_));
 sky130_fd_sc_hd__a32o_1 _12821_ (.A1(\cur_mb_mem[9][2] ),
    .A2(_06112_),
    .A3(_05910_),
    .B1(_06436_),
    .B2(\cur_mb_mem[158][2] ),
    .X(_07866_));
 sky130_fd_sc_hd__a32o_1 _12822_ (.A1(\cur_mb_mem[186][2] ),
    .A2(_05958_),
    .A3(_06036_),
    .B1(_06393_),
    .B2(\cur_mb_mem[34][2] ),
    .X(_07867_));
 sky130_fd_sc_hd__or4_2 _12823_ (.A(_07864_),
    .B(_07865_),
    .C(_07866_),
    .D(_07867_),
    .X(_07868_));
 sky130_fd_sc_hd__and3_1 _12824_ (.A(\cur_mb_mem[85][2] ),
    .B(_06927_),
    .C(_06794_),
    .X(_07869_));
 sky130_fd_sc_hd__and3_1 _12825_ (.A(\cur_mb_mem[171][2] ),
    .B(_06387_),
    .C(_07001_),
    .X(_07870_));
 sky130_fd_sc_hd__and3_1 _12826_ (.A(\cur_mb_mem[1][2] ),
    .B(_07096_),
    .C(_05993_),
    .X(_07871_));
 sky130_fd_sc_hd__a2111o_2 _12827_ (.A1(\cur_mb_mem[100][2] ),
    .A2(_06028_),
    .B1(_07869_),
    .C1(_07870_),
    .D1(_07871_),
    .X(_07872_));
 sky130_fd_sc_hd__and3_1 _12828_ (.A(\cur_mb_mem[116][2] ),
    .B(_06026_),
    .C(_06731_),
    .X(_07873_));
 sky130_fd_sc_hd__and3_2 _12829_ (.A(\cur_mb_mem[202][2] ),
    .B(_06442_),
    .C(_06986_),
    .X(_07874_));
 sky130_fd_sc_hd__and3_1 _12830_ (.A(\cur_mb_mem[252][2] ),
    .B(_06032_),
    .C(_06321_),
    .X(_07875_));
 sky130_fd_sc_hd__and3_1 _12831_ (.A(\cur_mb_mem[13][2] ),
    .B(_06300_),
    .C(_06011_),
    .X(_07876_));
 sky130_fd_sc_hd__or4_1 _12832_ (.A(_07873_),
    .B(_07874_),
    .C(_07875_),
    .D(_07876_),
    .X(_07877_));
 sky130_fd_sc_hd__and3_1 _12833_ (.A(\cur_mb_mem[181][2] ),
    .B(_06877_),
    .C(_06153_),
    .X(_07878_));
 sky130_fd_sc_hd__and3_1 _12834_ (.A(\cur_mb_mem[209][2] ),
    .B(_05947_),
    .C(_06251_),
    .X(_07879_));
 sky130_fd_sc_hd__and3_1 _12835_ (.A(\cur_mb_mem[200][2] ),
    .B(_06774_),
    .C(_06091_),
    .X(_07880_));
 sky130_fd_sc_hd__a2111o_4 _12836_ (.A1(\cur_mb_mem[14][2] ),
    .A2(_06367_),
    .B1(_07878_),
    .C1(_07879_),
    .D1(_07880_),
    .X(_07881_));
 sky130_fd_sc_hd__and3_1 _12837_ (.A(\cur_mb_mem[165][2] ),
    .B(_05922_),
    .C(_07279_),
    .X(_07882_));
 sky130_fd_sc_hd__and3_1 _12838_ (.A(\cur_mb_mem[126][2] ),
    .B(_07253_),
    .C(_07084_),
    .X(_07883_));
 sky130_fd_sc_hd__and3_1 _12839_ (.A(\cur_mb_mem[73][2] ),
    .B(_05893_),
    .C(_06023_),
    .X(_07884_));
 sky130_fd_sc_hd__a2111o_2 _12840_ (.A1(\cur_mb_mem[67][2] ),
    .A2(_06429_),
    .B1(_07882_),
    .C1(_07883_),
    .D1(_07884_),
    .X(_07885_));
 sky130_fd_sc_hd__or4_2 _12841_ (.A(_07872_),
    .B(_07877_),
    .C(_07881_),
    .D(_07885_),
    .X(_07886_));
 sky130_fd_sc_hd__a32o_1 _12842_ (.A1(\cur_mb_mem[204][2] ),
    .A2(_05938_),
    .A3(_06093_),
    .B1(_06383_),
    .B2(\cur_mb_mem[131][2] ),
    .X(_07887_));
 sky130_fd_sc_hd__a32o_1 _12843_ (.A1(\cur_mb_mem[54][2] ),
    .A2(_05057_),
    .A3(_06187_),
    .B1(_06088_),
    .B2(\cur_mb_mem[35][2] ),
    .X(_07888_));
 sky130_fd_sc_hd__nor2_1 _12844_ (.A(_07887_),
    .B(_07888_),
    .Y(_07889_));
 sky130_fd_sc_hd__a32o_2 _12845_ (.A1(\cur_mb_mem[113][2] ),
    .A2(_06053_),
    .A3(_05994_),
    .B1(_06402_),
    .B2(\cur_mb_mem[155][2] ),
    .X(_07890_));
 sky130_fd_sc_hd__a221oi_1 _12846_ (.A1(\cur_mb_mem[244][2] ),
    .A2(_06167_),
    .B1(_06290_),
    .B2(\cur_mb_mem[3][2] ),
    .C1(_07890_),
    .Y(_07891_));
 sky130_fd_sc_hd__or4bb_2 _12847_ (.A(_07868_),
    .B(_07886_),
    .C_N(_07889_),
    .D_N(_07891_),
    .X(_07892_));
 sky130_fd_sc_hd__or4_2 _12848_ (.A(_07853_),
    .B(_07854_),
    .C(_07863_),
    .D(_07892_),
    .X(_07893_));
 sky130_fd_sc_hd__a32o_1 _12849_ (.A1(\cur_mb_mem[247][2] ),
    .A2(_04431_),
    .A3(_06098_),
    .B1(_06248_),
    .B2(\cur_mb_mem[237][2] ),
    .X(_07894_));
 sky130_fd_sc_hd__a32o_1 _12850_ (.A1(\cur_mb_mem[175][2] ),
    .A2(_04424_),
    .A3(_06426_),
    .B1(_06447_),
    .B2(\cur_mb_mem[215][2] ),
    .X(_07895_));
 sky130_fd_sc_hd__a2111o_2 _12851_ (.A1(\cur_mb_mem[127][2] ),
    .A2(_06101_),
    .B1(_07894_),
    .C1(_07895_),
    .D1(_06185_),
    .X(_07896_));
 sky130_fd_sc_hd__a22o_1 _12852_ (.A1(\cur_mb_mem[242][2] ),
    .A2(_06335_),
    .B1(_06195_),
    .B2(\cur_mb_mem[164][2] ),
    .X(_07897_));
 sky130_fd_sc_hd__a221o_1 _12853_ (.A1(\cur_mb_mem[216][2] ),
    .A2(_06317_),
    .B1(_06433_),
    .B2(\cur_mb_mem[144][2] ),
    .C1(_07897_),
    .X(_07898_));
 sky130_fd_sc_hd__a22o_1 _12854_ (.A1(\cur_mb_mem[232][2] ),
    .A2(_06463_),
    .B1(_06117_),
    .B2(\cur_mb_mem[234][2] ),
    .X(_07899_));
 sky130_fd_sc_hd__a221o_1 _12855_ (.A1(\cur_mb_mem[15][2] ),
    .A2(_06295_),
    .B1(_06211_),
    .B2(\cur_mb_mem[134][2] ),
    .C1(_07899_),
    .X(_07900_));
 sky130_fd_sc_hd__a22o_1 _12856_ (.A1(\cur_mb_mem[226][2] ),
    .A2(_06256_),
    .B1(_06180_),
    .B2(\cur_mb_mem[231][2] ),
    .X(_07901_));
 sky130_fd_sc_hd__a32o_1 _12857_ (.A1(\cur_mb_mem[235][2] ),
    .A2(_06261_),
    .A3(_06224_),
    .B1(_06344_),
    .B2(\cur_mb_mem[37][2] ),
    .X(_07902_));
 sky130_fd_sc_hd__a32o_1 _12858_ (.A1(\cur_mb_mem[227][2] ),
    .A2(_06063_),
    .A3(_06224_),
    .B1(_06020_),
    .B2(\cur_mb_mem[177][2] ),
    .X(_07903_));
 sky130_fd_sc_hd__a22o_1 _12859_ (.A1(\cur_mb_mem[184][2] ),
    .A2(_06479_),
    .B1(_06160_),
    .B2(\cur_mb_mem[246][2] ),
    .X(_07904_));
 sky130_fd_sc_hd__or4_1 _12860_ (.A(_07901_),
    .B(_07902_),
    .C(_07903_),
    .D(_07904_),
    .X(_07905_));
 sky130_fd_sc_hd__and3_1 _12861_ (.A(\cur_mb_mem[172][2] ),
    .B(_06937_),
    .C(_07001_),
    .X(_07906_));
 sky130_fd_sc_hd__and3_1 _12862_ (.A(\cur_mb_mem[43][2] ),
    .B(_06942_),
    .C(_06044_),
    .X(_07907_));
 sky130_fd_sc_hd__and3_1 _12863_ (.A(\cur_mb_mem[88][2] ),
    .B(_06774_),
    .C(_07277_),
    .X(_07908_));
 sky130_fd_sc_hd__a2111o_1 _12864_ (.A1(\cur_mb_mem[61][2] ),
    .A2(_06359_),
    .B1(_07906_),
    .C1(_07907_),
    .D1(_07908_),
    .X(_07909_));
 sky130_fd_sc_hd__and3_2 _12865_ (.A(\cur_mb_mem[245][2] ),
    .B(_06902_),
    .C(_06153_),
    .X(_07910_));
 sky130_fd_sc_hd__and3_1 _12866_ (.A(\cur_mb_mem[112][2] ),
    .B(_07253_),
    .C(_06315_),
    .X(_07911_));
 sky130_fd_sc_hd__and3_1 _12867_ (.A(\cur_mb_mem[72][2] ),
    .B(_06774_),
    .C(_06023_),
    .X(_07912_));
 sky130_fd_sc_hd__a2111o_1 _12868_ (.A1(\cur_mb_mem[138][2] ),
    .A2(_05934_),
    .B1(_07910_),
    .C1(_07911_),
    .D1(_07912_),
    .X(_07913_));
 sky130_fd_sc_hd__and3_1 _12869_ (.A(\cur_mb_mem[133][2] ),
    .B(_06859_),
    .C(_06153_),
    .X(_07914_));
 sky130_fd_sc_hd__and3_1 _12870_ (.A(\cur_mb_mem[117][2] ),
    .B(_07253_),
    .C(_07279_),
    .X(_07915_));
 sky130_fd_sc_hd__and3_1 _12871_ (.A(\cur_mb_mem[120][2] ),
    .B(_06774_),
    .C(_07021_),
    .X(_07916_));
 sky130_fd_sc_hd__a2111o_1 _12872_ (.A1(\cur_mb_mem[97][2] ),
    .A2(_06077_),
    .B1(_07914_),
    .C1(_07915_),
    .D1(_07916_),
    .X(_07917_));
 sky130_fd_sc_hd__and3_1 _12873_ (.A(\cur_mb_mem[196][2] ),
    .B(_06166_),
    .C(_06352_),
    .X(_07918_));
 sky130_fd_sc_hd__and3_1 _12874_ (.A(\cur_mb_mem[198][2] ),
    .B(_06140_),
    .C(_06352_),
    .X(_07919_));
 sky130_fd_sc_hd__and3_1 _12875_ (.A(\cur_mb_mem[208][2] ),
    .B(_06814_),
    .C(_05970_),
    .X(_07920_));
 sky130_fd_sc_hd__and3_2 _12876_ (.A(\cur_mb_mem[75][2] ),
    .B(_06387_),
    .C(_06057_),
    .X(_07921_));
 sky130_fd_sc_hd__or4_2 _12877_ (.A(_07918_),
    .B(_07919_),
    .C(_07920_),
    .D(_07921_),
    .X(_07922_));
 sky130_fd_sc_hd__or4_4 _12878_ (.A(_07909_),
    .B(_07913_),
    .C(_07917_),
    .D(_07922_),
    .X(_07923_));
 sky130_fd_sc_hd__or4_2 _12879_ (.A(_07898_),
    .B(_07900_),
    .C(_07905_),
    .D(_07923_),
    .X(_07924_));
 sky130_fd_sc_hd__and3_1 _12880_ (.A(\cur_mb_mem[169][2] ),
    .B(_06723_),
    .C(_06755_),
    .X(_07925_));
 sky130_fd_sc_hd__and3_1 _12881_ (.A(\cur_mb_mem[168][2] ),
    .B(_06832_),
    .C(_06192_),
    .X(_07926_));
 sky130_fd_sc_hd__and3_1 _12882_ (.A(\cur_mb_mem[33][2] ),
    .B(_06044_),
    .C(_06251_),
    .X(_07927_));
 sky130_fd_sc_hd__a2111o_1 _12883_ (.A1(\cur_mb_mem[42][2] ),
    .A2(_06441_),
    .B1(_07925_),
    .C1(_07926_),
    .D1(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__and3_1 _12884_ (.A(\cur_mb_mem[102][2] ),
    .B(_06268_),
    .C(_06199_),
    .X(_07929_));
 sky130_fd_sc_hd__and3_1 _12885_ (.A(\cur_mb_mem[193][2] ),
    .B(_06967_),
    .C(_06912_),
    .X(_07930_));
 sky130_fd_sc_hd__and3_1 _12886_ (.A(\cur_mb_mem[96][2] ),
    .B(_06413_),
    .C(_06315_),
    .X(_07931_));
 sky130_fd_sc_hd__a2111o_1 _12887_ (.A1(\cur_mb_mem[74][2] ),
    .A2(_06417_),
    .B1(_07929_),
    .C1(_07930_),
    .D1(_07931_),
    .X(_07932_));
 sky130_fd_sc_hd__and3_2 _12888_ (.A(\cur_mb_mem[218][2] ),
    .B(_06960_),
    .C(_06150_),
    .X(_07933_));
 sky130_fd_sc_hd__and3_1 _12889_ (.A(\cur_mb_mem[137][2] ),
    .B(_06834_),
    .C(_06859_),
    .X(_07934_));
 sky130_fd_sc_hd__and3_1 _12890_ (.A(\cur_mb_mem[179][2] ),
    .B(_06086_),
    .C(_06216_),
    .X(_07935_));
 sky130_fd_sc_hd__a2111o_1 _12891_ (.A1(\cur_mb_mem[152][2] ),
    .A2(_06394_),
    .B1(_07933_),
    .C1(_07934_),
    .D1(_07935_),
    .X(_07936_));
 sky130_fd_sc_hd__and3_1 _12892_ (.A(\cur_mb_mem[109][2] ),
    .B(_06413_),
    .C(_06056_),
    .X(_07937_));
 sky130_fd_sc_hd__and3_1 _12893_ (.A(\cur_mb_mem[84][2] ),
    .B(_06215_),
    .C(_07277_),
    .X(_07938_));
 sky130_fd_sc_hd__and3_1 _12894_ (.A(\cur_mb_mem[251][2] ),
    .B(_07137_),
    .C(_05918_),
    .X(_07939_));
 sky130_fd_sc_hd__a2111o_1 _12895_ (.A1(\cur_mb_mem[110][2] ),
    .A2(_06047_),
    .B1(_07937_),
    .C1(_07938_),
    .D1(_07939_),
    .X(_07940_));
 sky130_fd_sc_hd__or4_4 _12896_ (.A(_07928_),
    .B(_07932_),
    .C(_07936_),
    .D(_07940_),
    .X(_07941_));
 sky130_fd_sc_hd__and3_1 _12897_ (.A(\cur_mb_mem[80][2] ),
    .B(_06230_),
    .C(_05970_),
    .X(_07942_));
 sky130_fd_sc_hd__and3_1 _12898_ (.A(\cur_mb_mem[17][2] ),
    .B(_06912_),
    .C(_06001_),
    .X(_07943_));
 sky130_fd_sc_hd__and3_1 _12899_ (.A(\cur_mb_mem[62][2] ),
    .B(_07235_),
    .C(_07084_),
    .X(_07944_));
 sky130_fd_sc_hd__a2111o_1 _12900_ (.A1(\cur_mb_mem[24][2] ),
    .A2(_06285_),
    .B1(_07942_),
    .C1(_07943_),
    .D1(_07944_),
    .X(_07945_));
 sky130_fd_sc_hd__and3_1 _12901_ (.A(\cur_mb_mem[130][2] ),
    .B(_06080_),
    .C(_06146_),
    .X(_07946_));
 sky130_fd_sc_hd__and3_2 _12902_ (.A(\cur_mb_mem[197][2] ),
    .B(_06967_),
    .C(_06794_),
    .X(_07947_));
 sky130_fd_sc_hd__and3_1 _12903_ (.A(\cur_mb_mem[92][2] ),
    .B(_06920_),
    .C(_06895_),
    .X(_07948_));
 sky130_fd_sc_hd__a2111o_1 _12904_ (.A1(\cur_mb_mem[161][2] ),
    .A2(_06334_),
    .B1(_07946_),
    .C1(_07947_),
    .D1(_07948_),
    .X(_07949_));
 sky130_fd_sc_hd__and3_1 _12905_ (.A(\cur_mb_mem[106][2] ),
    .B(_06960_),
    .C(_06268_),
    .X(_07950_));
 sky130_fd_sc_hd__and3_1 _12906_ (.A(\cur_mb_mem[188][2] ),
    .B(_06937_),
    .C(_06877_),
    .X(_07951_));
 sky130_fd_sc_hd__and3_1 _12907_ (.A(\cur_mb_mem[82][2] ),
    .B(_07099_),
    .C(_07277_),
    .X(_07952_));
 sky130_fd_sc_hd__a2111o_1 _12908_ (.A1(\cur_mb_mem[44][2] ),
    .A2(_06399_),
    .B1(_07950_),
    .C1(_07951_),
    .D1(_07952_),
    .X(_07953_));
 sky130_fd_sc_hd__and3_1 _12909_ (.A(\cur_mb_mem[254][2] ),
    .B(_06902_),
    .C(_07084_),
    .X(_07954_));
 sky130_fd_sc_hd__and3_1 _12910_ (.A(\cur_mb_mem[150][2] ),
    .B(_06191_),
    .C(_07100_),
    .X(_07955_));
 sky130_fd_sc_hd__and3_1 _12911_ (.A(\cur_mb_mem[212][2] ),
    .B(_05890_),
    .C(_05941_),
    .X(_07956_));
 sky130_fd_sc_hd__a2111o_4 _12912_ (.A1(\cur_mb_mem[253][2] ),
    .A2(_06034_),
    .B1(_07954_),
    .C1(_07955_),
    .D1(_07956_),
    .X(_07957_));
 sky130_fd_sc_hd__or4_2 _12913_ (.A(_07945_),
    .B(_07949_),
    .C(_07953_),
    .D(_07957_),
    .X(_07958_));
 sky130_fd_sc_hd__and3_1 _12914_ (.A(\cur_mb_mem[93][2] ),
    .B(_06008_),
    .C(_06033_),
    .X(_07959_));
 sky130_fd_sc_hd__and3_1 _12915_ (.A(\cur_mb_mem[220][2] ),
    .B(_06321_),
    .C(_06802_),
    .X(_07960_));
 sky130_fd_sc_hd__and3_1 _12916_ (.A(\cur_mb_mem[174][2] ),
    .B(_06366_),
    .C(_06333_),
    .X(_07961_));
 sky130_fd_sc_hd__and3_1 _12917_ (.A(\cur_mb_mem[206][2] ),
    .B(_06046_),
    .C(_06456_),
    .X(_07962_));
 sky130_fd_sc_hd__or4_1 _12918_ (.A(_07959_),
    .B(_07960_),
    .C(_07961_),
    .D(_07962_),
    .X(_07963_));
 sky130_fd_sc_hd__and3_1 _12919_ (.A(\cur_mb_mem[32][2] ),
    .B(_06952_),
    .C(_06772_),
    .X(_07964_));
 sky130_fd_sc_hd__and3_1 _12920_ (.A(\cur_mb_mem[8][2] ),
    .B(_07096_),
    .C(_06832_),
    .X(_07965_));
 sky130_fd_sc_hd__and3_1 _12921_ (.A(\cur_mb_mem[156][2] ),
    .B(_06920_),
    .C(_07100_),
    .X(_07966_));
 sky130_fd_sc_hd__a2111o_1 _12922_ (.A1(\cur_mb_mem[211][2] ),
    .A2(_06349_),
    .B1(_07964_),
    .C1(_07965_),
    .D1(_07966_),
    .X(_07967_));
 sky130_fd_sc_hd__and3_1 _12923_ (.A(\cur_mb_mem[157][2] ),
    .B(_06056_),
    .C(_06152_),
    .X(_07968_));
 sky130_fd_sc_hd__and3_1 _12924_ (.A(\cur_mb_mem[21][2] ),
    .B(_06001_),
    .C(_06153_),
    .X(_07969_));
 sky130_fd_sc_hd__and3_1 _12925_ (.A(\cur_mb_mem[249][2] ),
    .B(_07137_),
    .C(_05893_),
    .X(_07970_));
 sky130_fd_sc_hd__a2111o_1 _12926_ (.A1(\cur_mb_mem[250][2] ),
    .A2(_06443_),
    .B1(_07968_),
    .C1(_07969_),
    .D1(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__and3_1 _12927_ (.A(\cur_mb_mem[213][2] ),
    .B(_05947_),
    .C(_07279_),
    .X(_07972_));
 sky130_fd_sc_hd__and3_1 _12928_ (.A(\cur_mb_mem[149][2] ),
    .B(_07100_),
    .C(_07279_),
    .X(_07973_));
 sky130_fd_sc_hd__and3_1 _12929_ (.A(\cur_mb_mem[107][2] ),
    .B(_05918_),
    .C(_06413_),
    .X(_07974_));
 sky130_fd_sc_hd__a2111o_1 _12930_ (.A1(\cur_mb_mem[6][2] ),
    .A2(_06203_),
    .B1(_07972_),
    .C1(_07973_),
    .D1(_07974_),
    .X(_07975_));
 sky130_fd_sc_hd__or4_4 _12931_ (.A(_07963_),
    .B(_07967_),
    .C(_07971_),
    .D(_07975_),
    .X(_07976_));
 sky130_fd_sc_hd__and3_1 _12932_ (.A(\cur_mb_mem[243][2] ),
    .B(_06902_),
    .C(_06086_),
    .X(_07977_));
 sky130_fd_sc_hd__and3_1 _12933_ (.A(\cur_mb_mem[229][2] ),
    .B(_07279_),
    .C(_06775_),
    .X(_07978_));
 sky130_fd_sc_hd__and3_1 _12934_ (.A(\cur_mb_mem[60][2] ),
    .B(_05056_),
    .C(_06920_),
    .X(_07979_));
 sky130_fd_sc_hd__a2111o_2 _12935_ (.A1(\cur_mb_mem[53][2] ),
    .A2(_06221_),
    .B1(_07977_),
    .C1(_07978_),
    .D1(_07979_),
    .X(_07980_));
 sky130_fd_sc_hd__and3_1 _12936_ (.A(\cur_mb_mem[207][2] ),
    .B(_04423_),
    .C(_06997_),
    .X(_07981_));
 sky130_fd_sc_hd__and3_1 _12937_ (.A(\cur_mb_mem[236][2] ),
    .B(_06920_),
    .C(_06775_),
    .X(_07982_));
 sky130_fd_sc_hd__and3_1 _12938_ (.A(\cur_mb_mem[167][2] ),
    .B(_05922_),
    .C(_06096_),
    .X(_07983_));
 sky130_fd_sc_hd__a2111o_1 _12939_ (.A1(\cur_mb_mem[79][2] ),
    .A2(_06122_),
    .B1(_07981_),
    .C1(_07982_),
    .D1(_07983_),
    .X(_07984_));
 sky130_fd_sc_hd__and3_1 _12940_ (.A(\cur_mb_mem[48][2] ),
    .B(_07235_),
    .C(_06315_),
    .X(_07985_));
 sky130_fd_sc_hd__and3_1 _12941_ (.A(\cur_mb_mem[241][2] ),
    .B(_07137_),
    .C(_05993_),
    .X(_07986_));
 sky130_fd_sc_hd__and3_1 _12942_ (.A(\cur_mb_mem[41][2] ),
    .B(_05893_),
    .C(_06044_),
    .X(_07987_));
 sky130_fd_sc_hd__a2111o_1 _12943_ (.A1(\cur_mb_mem[182][2] ),
    .A2(_06205_),
    .B1(_07985_),
    .C1(_07986_),
    .D1(_07987_),
    .X(_07988_));
 sky130_fd_sc_hd__and3_1 _12944_ (.A(\cur_mb_mem[26][2] ),
    .B(_05957_),
    .C(_06235_),
    .X(_07989_));
 sky130_fd_sc_hd__and3_1 _12945_ (.A(\cur_mb_mem[240][2] ),
    .B(_06165_),
    .C(_05970_),
    .X(_07990_));
 sky130_fd_sc_hd__and3_1 _12946_ (.A(\cur_mb_mem[183][2] ),
    .B(_06760_),
    .C(_06372_),
    .X(_07991_));
 sky130_fd_sc_hd__and3_1 _12947_ (.A(\cur_mb_mem[23][2] ),
    .B(_06896_),
    .C(_06001_),
    .X(_07992_));
 sky130_fd_sc_hd__or4_1 _12948_ (.A(_07989_),
    .B(_07990_),
    .C(_07991_),
    .D(_07992_),
    .X(_07993_));
 sky130_fd_sc_hd__or4_2 _12949_ (.A(_07980_),
    .B(_07984_),
    .C(_07988_),
    .D(_07993_),
    .X(_07994_));
 sky130_fd_sc_hd__or4_1 _12950_ (.A(_07941_),
    .B(_07958_),
    .C(_07976_),
    .D(_07994_),
    .X(_07995_));
 sky130_fd_sc_hd__and3_1 _12951_ (.A(\cur_mb_mem[63][2] ),
    .B(_06149_),
    .C(_06198_),
    .X(_07996_));
 sky130_fd_sc_hd__and3_1 _12952_ (.A(\cur_mb_mem[224][2] ),
    .B(_06748_),
    .C(_06775_),
    .X(_07997_));
 sky130_fd_sc_hd__and3_1 _12953_ (.A(\cur_mb_mem[191][2] ),
    .B(_04423_),
    .C(_06216_),
    .X(_07998_));
 sky130_fd_sc_hd__a2111o_4 _12954_ (.A1(\cur_mb_mem[255][2] ),
    .A2(_06304_),
    .B1(_07996_),
    .C1(_07997_),
    .D1(_07998_),
    .X(_07999_));
 sky130_fd_sc_hd__and3_1 _12955_ (.A(\cur_mb_mem[111][2] ),
    .B(_06068_),
    .C(_06027_),
    .X(_08000_));
 sky130_fd_sc_hd__and3_1 _12956_ (.A(\cur_mb_mem[71][2] ),
    .B(_06428_),
    .C(_06461_),
    .X(_08001_));
 sky130_fd_sc_hd__and3_1 _12957_ (.A(\cur_mb_mem[103][2] ),
    .B(_06313_),
    .C(_06461_),
    .X(_08002_));
 sky130_fd_sc_hd__and3_1 _12958_ (.A(\cur_mb_mem[47][2] ),
    .B(_06466_),
    .C(_06343_),
    .X(_08003_));
 sky130_fd_sc_hd__or4_4 _12959_ (.A(_08000_),
    .B(_08001_),
    .C(_08002_),
    .D(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__and3_1 _12960_ (.A(\cur_mb_mem[40][2] ),
    .B(_06832_),
    .C(_06087_),
    .X(_08005_));
 sky130_fd_sc_hd__and3_1 _12961_ (.A(\cur_mb_mem[98][2] ),
    .B(_07099_),
    .C(_06413_),
    .X(_08006_));
 sky130_fd_sc_hd__and3_1 _12962_ (.A(\cur_mb_mem[210][2] ),
    .B(_07099_),
    .C(_05941_),
    .X(_08007_));
 sky130_fd_sc_hd__a2111o_1 _12963_ (.A1(\cur_mb_mem[91][2] ),
    .A2(_06361_),
    .B1(_08005_),
    .C1(_08006_),
    .D1(_08007_),
    .X(_08008_));
 sky130_fd_sc_hd__and3_2 _12964_ (.A(\cur_mb_mem[238][2] ),
    .B(_07084_),
    .C(_06065_),
    .X(_08009_));
 sky130_fd_sc_hd__and3_1 _12965_ (.A(\cur_mb_mem[151][2] ),
    .B(_05978_),
    .C(_06096_),
    .X(_08010_));
 sky130_fd_sc_hd__and3_1 _12966_ (.A(\cur_mb_mem[123][2] ),
    .B(_05918_),
    .C(_07021_),
    .X(_08011_));
 sky130_fd_sc_hd__a2111o_1 _12967_ (.A1(\cur_mb_mem[68][2] ),
    .A2(_06234_),
    .B1(_08009_),
    .C1(_08010_),
    .D1(_08011_),
    .X(_08012_));
 sky130_fd_sc_hd__or4_4 _12968_ (.A(_07999_),
    .B(_08004_),
    .C(_08008_),
    .D(_08012_),
    .X(_08013_));
 sky130_fd_sc_hd__and3_2 _12969_ (.A(\cur_mb_mem[146][2] ),
    .B(_06908_),
    .C(_06152_),
    .X(_08014_));
 sky130_fd_sc_hd__and3_1 _12970_ (.A(\cur_mb_mem[199][2] ),
    .B(_06997_),
    .C(_07195_),
    .X(_08015_));
 sky130_fd_sc_hd__and3_1 _12971_ (.A(\cur_mb_mem[87][2] ),
    .B(_07277_),
    .C(_06096_),
    .X(_08016_));
 sky130_fd_sc_hd__a2111o_1 _12972_ (.A1(\cur_mb_mem[135][2] ),
    .A2(_06462_),
    .B1(_08014_),
    .C1(_08015_),
    .D1(_08016_),
    .X(_08017_));
 sky130_fd_sc_hd__and3_1 _12973_ (.A(\cur_mb_mem[76][2] ),
    .B(_06937_),
    .C(_06057_),
    .X(_08018_));
 sky130_fd_sc_hd__and3_4 _12974_ (.A(\cur_mb_mem[114][2] ),
    .B(_06380_),
    .C(_07253_),
    .X(_08019_));
 sky130_fd_sc_hd__and3_1 _12975_ (.A(\cur_mb_mem[49][2] ),
    .B(_05056_),
    .C(_05993_),
    .X(_08020_));
 sky130_fd_sc_hd__a2111o_1 _12976_ (.A1(\cur_mb_mem[225][2] ),
    .A2(_05998_),
    .B1(_08018_),
    .C1(_08019_),
    .D1(_08020_),
    .X(_08021_));
 sky130_fd_sc_hd__and3_1 _12977_ (.A(\cur_mb_mem[7][2] ),
    .B(_07096_),
    .C(_07195_),
    .X(_08022_));
 sky130_fd_sc_hd__and3_1 _12978_ (.A(\cur_mb_mem[119][2] ),
    .B(_07253_),
    .C(_07195_),
    .X(_08023_));
 sky130_fd_sc_hd__and3_1 _12979_ (.A(\cur_mb_mem[233][2] ),
    .B(_05893_),
    .C(_06065_),
    .X(_08024_));
 sky130_fd_sc_hd__a2111o_1 _12980_ (.A1(\cur_mb_mem[248][2] ),
    .A2(_06411_),
    .B1(_08022_),
    .C1(_08023_),
    .D1(_08024_),
    .X(_08025_));
 sky130_fd_sc_hd__and3_1 _12981_ (.A(\cur_mb_mem[55][2] ),
    .B(_05056_),
    .C(_06096_),
    .X(_08026_));
 sky130_fd_sc_hd__and3_1 _12982_ (.A(\cur_mb_mem[143][2] ),
    .B(_04423_),
    .C(_05935_),
    .X(_08027_));
 sky130_fd_sc_hd__and3_1 _12983_ (.A(\cur_mb_mem[228][2] ),
    .B(_05890_),
    .C(_06065_),
    .X(_08028_));
 sky130_fd_sc_hd__a2111o_1 _12984_ (.A1(\cur_mb_mem[39][2] ),
    .A2(_06373_),
    .B1(_08026_),
    .C1(_08027_),
    .D1(_08028_),
    .X(_08029_));
 sky130_fd_sc_hd__or4_1 _12985_ (.A(_08017_),
    .B(_08021_),
    .C(_08025_),
    .D(_08029_),
    .X(_08030_));
 sky130_fd_sc_hd__and3_1 _12986_ (.A(\cur_mb_mem[173][2] ),
    .B(_06246_),
    .C(_07001_),
    .X(_08031_));
 sky130_fd_sc_hd__and3_1 _12987_ (.A(\cur_mb_mem[205][2] ),
    .B(_06246_),
    .C(_06997_),
    .X(_08032_));
 sky130_fd_sc_hd__and3_1 _12988_ (.A(\cur_mb_mem[139][2] ),
    .B(_05918_),
    .C(_05935_),
    .X(_08033_));
 sky130_fd_sc_hd__a2111o_2 _12989_ (.A1(\cur_mb_mem[142][2] ),
    .A2(_06487_),
    .B1(_08031_),
    .C1(_08032_),
    .D1(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__and3_1 _12990_ (.A(\cur_mb_mem[162][2] ),
    .B(_06380_),
    .C(_07001_),
    .X(_08035_));
 sky130_fd_sc_hd__and3_1 _12991_ (.A(\cur_mb_mem[239][2] ),
    .B(_04423_),
    .C(_06775_),
    .X(_08036_));
 sky130_fd_sc_hd__and3_1 _12992_ (.A(\cur_mb_mem[230][2] ),
    .B(_06186_),
    .C(_06065_),
    .X(_08037_));
 sky130_fd_sc_hd__a2111o_1 _12993_ (.A1(\cur_mb_mem[56][2] ),
    .A2(_06351_),
    .B1(_08035_),
    .C1(_08036_),
    .D1(_08037_),
    .X(_08038_));
 sky130_fd_sc_hd__and3_1 _12994_ (.A(\cur_mb_mem[94][2] ),
    .B(_07277_),
    .C(_07084_),
    .X(_08039_));
 sky130_fd_sc_hd__and3_1 _12995_ (.A(\cur_mb_mem[187][2] ),
    .B(_05918_),
    .C(_06216_),
    .X(_08040_));
 sky130_fd_sc_hd__and3_1 _12996_ (.A(\cur_mb_mem[189][2] ),
    .B(_05945_),
    .C(_06036_),
    .X(_08041_));
 sky130_fd_sc_hd__a2111o_1 _12997_ (.A1(\cur_mb_mem[118][2] ),
    .A2(_06141_),
    .B1(_08039_),
    .C1(_08040_),
    .D1(_08041_),
    .X(_08042_));
 sky130_fd_sc_hd__and3_1 _12998_ (.A(\cur_mb_mem[59][2] ),
    .B(_05056_),
    .C(_05918_),
    .X(_08043_));
 sky130_fd_sc_hd__and3_1 _12999_ (.A(\cur_mb_mem[195][2] ),
    .B(_06062_),
    .C(_06091_),
    .X(_08044_));
 sky130_fd_sc_hd__and3_1 _13000_ (.A(\cur_mb_mem[99][2] ),
    .B(_06298_),
    .C(_06062_),
    .X(_08045_));
 sky130_fd_sc_hd__a2111o_1 _13001_ (.A1(\cur_mb_mem[50][2] ),
    .A2(_06172_),
    .B1(_08043_),
    .C1(_08044_),
    .D1(_08045_),
    .X(_08046_));
 sky130_fd_sc_hd__or4_2 _13002_ (.A(_08034_),
    .B(_08038_),
    .C(_08042_),
    .D(_08046_),
    .X(_08047_));
 sky130_fd_sc_hd__and3_1 _13003_ (.A(\cur_mb_mem[66][2] ),
    .B(_07099_),
    .C(_06023_),
    .X(_08048_));
 sky130_fd_sc_hd__and3_1 _13004_ (.A(\cur_mb_mem[90][2] ),
    .B(_05905_),
    .C(_07277_),
    .X(_08049_));
 sky130_fd_sc_hd__and3_1 _13005_ (.A(\cur_mb_mem[163][2] ),
    .B(_06062_),
    .C(_05922_),
    .X(_08050_));
 sky130_fd_sc_hd__a2111o_1 _13006_ (.A1(\cur_mb_mem[83][2] ),
    .A2(_06379_),
    .B1(_08048_),
    .C1(_08049_),
    .D1(_08050_),
    .X(_08051_));
 sky130_fd_sc_hd__and3_1 _13007_ (.A(\cur_mb_mem[2][2] ),
    .B(_07096_),
    .C(_07099_),
    .X(_08052_));
 sky130_fd_sc_hd__and3_1 _13008_ (.A(\cur_mb_mem[115][2] ),
    .B(_06086_),
    .C(_07021_),
    .X(_08053_));
 sky130_fd_sc_hd__and3_1 _13009_ (.A(\cur_mb_mem[147][2] ),
    .B(_06062_),
    .C(_05978_),
    .X(_08054_));
 sky130_fd_sc_hd__a2111o_1 _13010_ (.A1(\cur_mb_mem[52][2] ),
    .A2(_06241_),
    .B1(_08052_),
    .C1(_08053_),
    .D1(_08054_),
    .X(_08055_));
 sky130_fd_sc_hd__and3_1 _13011_ (.A(\cur_mb_mem[121][2] ),
    .B(_05893_),
    .C(_07021_),
    .X(_08056_));
 sky130_fd_sc_hd__and3_1 _13012_ (.A(\cur_mb_mem[140][2] ),
    .B(_05937_),
    .C(_05935_),
    .X(_08057_));
 sky130_fd_sc_hd__and3_1 _13013_ (.A(\cur_mb_mem[178][2] ),
    .B(_06283_),
    .C(_06036_),
    .X(_08058_));
 sky130_fd_sc_hd__a2111o_1 _13014_ (.A1(\cur_mb_mem[104][2] ),
    .A2(_05985_),
    .B1(_08056_),
    .C1(_08057_),
    .D1(_08058_),
    .X(_08059_));
 sky130_fd_sc_hd__and3_1 _13015_ (.A(\cur_mb_mem[18][2] ),
    .B(_07099_),
    .C(_05975_),
    .X(_08060_));
 sky130_fd_sc_hd__and3_1 _13016_ (.A(\cur_mb_mem[5][2] ),
    .B(_06112_),
    .C(_07279_),
    .X(_08061_));
 sky130_fd_sc_hd__and3_1 _13017_ (.A(\cur_mb_mem[153][2] ),
    .B(_05910_),
    .C(_05978_),
    .X(_08062_));
 sky130_fd_sc_hd__a2111o_1 _13018_ (.A1(\cur_mb_mem[30][2] ),
    .A2(_06002_),
    .B1(_08060_),
    .C1(_08061_),
    .D1(_08062_),
    .X(_08063_));
 sky130_fd_sc_hd__or4_4 _13019_ (.A(_08051_),
    .B(_08055_),
    .C(_08059_),
    .D(_08063_),
    .X(_08064_));
 sky130_fd_sc_hd__or4_1 _13020_ (.A(_08013_),
    .B(_08030_),
    .C(_08047_),
    .D(_08064_),
    .X(_08065_));
 sky130_fd_sc_hd__or4_4 _13021_ (.A(_07896_),
    .B(_07924_),
    .C(_07995_),
    .D(_08065_),
    .X(_08066_));
 sky130_fd_sc_hd__nor4_1 _13022_ (.A(_07837_),
    .B(_07852_),
    .C(_07893_),
    .D(_08066_),
    .Y(_08067_));
 sky130_fd_sc_hd__nor3_2 _13023_ (.A(net99),
    .B(_07820_),
    .C(net211),
    .Y(_08068_));
 sky130_fd_sc_hd__o21a_1 _13024_ (.A1(_07820_),
    .A2(net211),
    .B1(net99),
    .X(_08069_));
 sky130_fd_sc_hd__a2111o_1 _13025_ (.A1(_07552_),
    .A2(_07553_),
    .B1(_07819_),
    .C1(_08068_),
    .D1(_08069_),
    .X(_08070_));
 sky130_fd_sc_hd__nand2_1 _13026_ (.A(net100),
    .B(_07818_),
    .Y(_08071_));
 sky130_fd_sc_hd__nor2_1 _13027_ (.A(net100),
    .B(_07818_),
    .Y(_08072_));
 sky130_fd_sc_hd__a21oi_1 _13028_ (.A1(_08071_),
    .A2(_08068_),
    .B1(_08072_),
    .Y(_08073_));
 sky130_fd_sc_hd__xor2_1 _13029_ (.A(net102),
    .B(_07009_),
    .X(_08074_));
 sky130_fd_sc_hd__a32o_1 _13030_ (.A1(\cur_mb_mem[123][4] ),
    .A2(_05919_),
    .A3(_06053_),
    .B1(_06394_),
    .B2(\cur_mb_mem[152][4] ),
    .X(_08075_));
 sky130_fd_sc_hd__and3_1 _13031_ (.A(\cur_mb_mem[125][4] ),
    .B(_05945_),
    .C(_06052_),
    .X(_08076_));
 sky130_fd_sc_hd__a31o_1 _13032_ (.A1(\cur_mb_mem[124][4] ),
    .A2(_05937_),
    .A3(_06118_),
    .B1(_08076_),
    .X(_08077_));
 sky130_fd_sc_hd__a32o_1 _13033_ (.A1(\cur_mb_mem[122][4] ),
    .A2(_05958_),
    .A3(_06118_),
    .B1(_06196_),
    .B2(\cur_mb_mem[132][4] ),
    .X(_08078_));
 sky130_fd_sc_hd__a211o_1 _13034_ (.A1(\cur_mb_mem[158][4] ),
    .A2(_06436_),
    .B1(_08077_),
    .C1(_08078_),
    .X(_08079_));
 sky130_fd_sc_hd__a211o_1 _13035_ (.A1(\cur_mb_mem[133][4] ),
    .A2(_06148_),
    .B1(_08075_),
    .C1(_08079_),
    .X(_08080_));
 sky130_fd_sc_hd__a32o_1 _13036_ (.A1(\cur_mb_mem[121][4] ),
    .A2(_06336_),
    .A3(_06053_),
    .B1(_06439_),
    .B2(\cur_mb_mem[112][4] ),
    .X(_08081_));
 sky130_fd_sc_hd__a221o_1 _13037_ (.A1(\cur_mb_mem[146][4] ),
    .A2(_06381_),
    .B1(_06231_),
    .B2(\cur_mb_mem[85][4] ),
    .C1(_08081_),
    .X(_08082_));
 sky130_fd_sc_hd__a22o_1 _13038_ (.A1(\cur_mb_mem[118][4] ),
    .A2(_06141_),
    .B1(_06209_),
    .B2(\cur_mb_mem[117][4] ),
    .X(_08083_));
 sky130_fd_sc_hd__a221o_1 _13039_ (.A1(\cur_mb_mem[116][4] ),
    .A2(_06239_),
    .B1(_06402_),
    .B2(\cur_mb_mem[155][4] ),
    .C1(_08083_),
    .X(_08084_));
 sky130_fd_sc_hd__or4_4 _13040_ (.A(_06185_),
    .B(_08080_),
    .C(_08082_),
    .D(_08084_),
    .X(_08085_));
 sky130_fd_sc_hd__and3_1 _13041_ (.A(\cur_mb_mem[16][4] ),
    .B(_06074_),
    .C(net232),
    .X(_08086_));
 sky130_fd_sc_hd__and3_1 _13042_ (.A(\cur_mb_mem[78][4] ),
    .B(_06428_),
    .C(_06366_),
    .X(_08087_));
 sky130_fd_sc_hd__and3_1 _13043_ (.A(\cur_mb_mem[18][4] ),
    .B(_06341_),
    .C(_06488_),
    .X(_08088_));
 sky130_fd_sc_hd__a2111o_1 _13044_ (.A1(\cur_mb_mem[17][4] ),
    .A2(_06318_),
    .B1(_08086_),
    .C1(_08087_),
    .D1(_08088_),
    .X(_08089_));
 sky130_fd_sc_hd__and3_1 _13045_ (.A(\cur_mb_mem[5][4] ),
    .B(_06365_),
    .C(_06131_),
    .X(_08090_));
 sky130_fd_sc_hd__and3_4 _13046_ (.A(\cur_mb_mem[190][4] ),
    .B(_06013_),
    .C(_06366_),
    .X(_08091_));
 sky130_fd_sc_hd__and3_1 _13047_ (.A(\cur_mb_mem[23][4] ),
    .B(_06461_),
    .C(_06475_),
    .X(_08092_));
 sky130_fd_sc_hd__a2111o_1 _13048_ (.A1(\cur_mb_mem[164][4] ),
    .A2(_06195_),
    .B1(_08090_),
    .C1(_08091_),
    .D1(_08092_),
    .X(_08093_));
 sky130_fd_sc_hd__and3_1 _13049_ (.A(\cur_mb_mem[29][4] ),
    .B(_06033_),
    .C(_06403_),
    .X(_08094_));
 sky130_fd_sc_hd__and3_1 _13050_ (.A(\cur_mb_mem[27][4] ),
    .B(_06003_),
    .C(_06488_),
    .X(_08095_));
 sky130_fd_sc_hd__and3_1 _13051_ (.A(\cur_mb_mem[1][4] ),
    .B(_06300_),
    .C(_06353_),
    .X(_08096_));
 sky130_fd_sc_hd__a2111o_1 _13052_ (.A1(\cur_mb_mem[19][4] ),
    .A2(_06282_),
    .B1(_08094_),
    .C1(_08095_),
    .D1(_08096_),
    .X(_08097_));
 sky130_fd_sc_hd__and3_1 _13053_ (.A(\cur_mb_mem[28][4] ),
    .B(_06422_),
    .C(_06488_),
    .X(_08098_));
 sky130_fd_sc_hd__and3_1 _13054_ (.A(\cur_mb_mem[4][4] ),
    .B(_06744_),
    .C(_06300_),
    .X(_08099_));
 sky130_fd_sc_hd__and3_1 _13055_ (.A(\cur_mb_mem[7][4] ),
    .B(_06707_),
    .C(_06372_),
    .X(_08100_));
 sky130_fd_sc_hd__a2111o_1 _13056_ (.A1(\cur_mb_mem[12][4] ),
    .A2(_05928_),
    .B1(_08098_),
    .C1(_08099_),
    .D1(_08100_),
    .X(_08101_));
 sky130_fd_sc_hd__or4_4 _13057_ (.A(_08089_),
    .B(_08093_),
    .C(_08097_),
    .D(_08101_),
    .X(_08102_));
 sky130_fd_sc_hd__and3_1 _13058_ (.A(\cur_mb_mem[3][4] ),
    .B(_06365_),
    .C(_06061_),
    .X(_08103_));
 sky130_fd_sc_hd__and3_1 _13059_ (.A(\cur_mb_mem[30][4] ),
    .B(_06366_),
    .C(_06403_),
    .X(_08104_));
 sky130_fd_sc_hd__and3_1 _13060_ (.A(\cur_mb_mem[24][4] ),
    .B(_05895_),
    .C(_06475_),
    .X(_08105_));
 sky130_fd_sc_hd__a2111o_1 _13061_ (.A1(\cur_mb_mem[26][4] ),
    .A2(_06449_),
    .B1(_08103_),
    .C1(_08104_),
    .D1(_08105_),
    .X(_08106_));
 sky130_fd_sc_hd__and3_1 _13062_ (.A(\cur_mb_mem[77][4] ),
    .B(_06033_),
    .C(_06428_),
    .X(_08107_));
 sky130_fd_sc_hd__and3_1 _13063_ (.A(\cur_mb_mem[66][4] ),
    .B(_06171_),
    .C(_06428_),
    .X(_08108_));
 sky130_fd_sc_hd__and3_1 _13064_ (.A(\cur_mb_mem[76][4] ),
    .B(_06718_),
    .C(_06121_),
    .X(_08109_));
 sky130_fd_sc_hd__a2111o_1 _13065_ (.A1(\cur_mb_mem[72][4] ),
    .A2(_06288_),
    .B1(_08107_),
    .C1(_08108_),
    .D1(_08109_),
    .X(_08110_));
 sky130_fd_sc_hd__and3_1 _13066_ (.A(\cur_mb_mem[22][4] ),
    .B(_06159_),
    .C(_06403_),
    .X(_08111_));
 sky130_fd_sc_hd__and3_1 _13067_ (.A(\cur_mb_mem[75][4] ),
    .B(_06003_),
    .C(_06143_),
    .X(_08112_));
 sky130_fd_sc_hd__and3_1 _13068_ (.A(\cur_mb_mem[9][4] ),
    .B(_06300_),
    .C(_06327_),
    .X(_08113_));
 sky130_fd_sc_hd__a2111o_1 _13069_ (.A1(\cur_mb_mem[14][4] ),
    .A2(_06367_),
    .B1(_08111_),
    .C1(_08112_),
    .D1(_08113_),
    .X(_08114_));
 sky130_fd_sc_hd__and3_1 _13070_ (.A(\cur_mb_mem[25][4] ),
    .B(_06038_),
    .C(_06488_),
    .X(_08115_));
 sky130_fd_sc_hd__and3_1 _13071_ (.A(\cur_mb_mem[2][4] ),
    .B(_06300_),
    .C(_06341_),
    .X(_08116_));
 sky130_fd_sc_hd__and3_1 _13072_ (.A(\cur_mb_mem[8][4] ),
    .B(_06707_),
    .C(_06478_),
    .X(_08117_));
 sky130_fd_sc_hd__a2111o_1 _13073_ (.A1(\cur_mb_mem[67][4] ),
    .A2(_06429_),
    .B1(_08115_),
    .C1(_08116_),
    .D1(_08117_),
    .X(_08118_));
 sky130_fd_sc_hd__or4_4 _13074_ (.A(_08106_),
    .B(_08110_),
    .C(_08114_),
    .D(_08118_),
    .X(_08119_));
 sky130_fd_sc_hd__and3_1 _13075_ (.A(\cur_mb_mem[113][4] ),
    .B(_06731_),
    .C(_06076_),
    .X(_08120_));
 sky130_fd_sc_hd__and3_1 _13076_ (.A(\cur_mb_mem[114][4] ),
    .B(_06171_),
    .C(_06731_),
    .X(_08121_));
 sky130_fd_sc_hd__and3_1 _13077_ (.A(\cur_mb_mem[119][4] ),
    .B(_06051_),
    .C(_06179_),
    .X(_08122_));
 sky130_fd_sc_hd__a2111o_1 _13078_ (.A1(\cur_mb_mem[43][4] ),
    .A2(_06006_),
    .B1(_08120_),
    .C1(_08121_),
    .D1(_08122_),
    .X(_08123_));
 sky130_fd_sc_hd__and3_1 _13079_ (.A(\cur_mb_mem[147][4] ),
    .B(_06061_),
    .C(_06188_),
    .X(_08124_));
 sky130_fd_sc_hd__and3_1 _13080_ (.A(\cur_mb_mem[126][4] ),
    .B(_06731_),
    .C(_06046_),
    .X(_08125_));
 sky130_fd_sc_hd__and3_1 _13081_ (.A(\cur_mb_mem[151][4] ),
    .B(_06434_),
    .C(_06179_),
    .X(_08126_));
 sky130_fd_sc_hd__a2111o_1 _13082_ (.A1(\cur_mb_mem[41][4] ),
    .A2(_06031_),
    .B1(_08124_),
    .C1(_08125_),
    .D1(_08126_),
    .X(_08127_));
 sky130_fd_sc_hd__and3_1 _13083_ (.A(\cur_mb_mem[156][4] ),
    .B(_06321_),
    .C(_06188_),
    .X(_08128_));
 sky130_fd_sc_hd__and3_1 _13084_ (.A(\cur_mb_mem[115][4] ),
    .B(_06355_),
    .C(_06051_),
    .X(_08129_));
 sky130_fd_sc_hd__and3_1 _13085_ (.A(\cur_mb_mem[120][4] ),
    .B(_06455_),
    .C(_06138_),
    .X(_08130_));
 sky130_fd_sc_hd__a2111o_1 _13086_ (.A1(\cur_mb_mem[150][4] ),
    .A2(_06189_),
    .B1(_08128_),
    .C1(_08129_),
    .D1(_08130_),
    .X(_08131_));
 sky130_fd_sc_hd__and3_2 _13087_ (.A(\cur_mb_mem[84][4] ),
    .B(_06744_),
    .C(_06378_),
    .X(_08132_));
 sky130_fd_sc_hd__and3_1 _13088_ (.A(\cur_mb_mem[149][4] ),
    .B(_06434_),
    .C(_06812_),
    .X(_08133_));
 sky130_fd_sc_hd__and3_1 _13089_ (.A(\cur_mb_mem[144][4] ),
    .B(_06747_),
    .C(_06772_),
    .X(_08134_));
 sky130_fd_sc_hd__a2111o_1 _13090_ (.A1(\cur_mb_mem[42][4] ),
    .A2(_06441_),
    .B1(_08132_),
    .C1(_08133_),
    .D1(_08134_),
    .X(_08135_));
 sky130_fd_sc_hd__or4_4 _13091_ (.A(_08123_),
    .B(_08127_),
    .C(_08131_),
    .D(_08135_),
    .X(_08136_));
 sky130_fd_sc_hd__and3_1 _13092_ (.A(\cur_mb_mem[179][4] ),
    .B(_06347_),
    .C(_06039_),
    .X(_08137_));
 sky130_fd_sc_hd__and3_1 _13093_ (.A(\cur_mb_mem[188][4] ),
    .B(_06718_),
    .C(_06039_),
    .X(_08138_));
 sky130_fd_sc_hd__and3_1 _13094_ (.A(\cur_mb_mem[172][4] ),
    .B(_06754_),
    .C(_06755_),
    .X(_08139_));
 sky130_fd_sc_hd__a2111o_1 _13095_ (.A1(\cur_mb_mem[189][4] ),
    .A2(_06014_),
    .B1(_08137_),
    .C1(_08138_),
    .D1(_08139_),
    .X(_08140_));
 sky130_fd_sc_hd__and3_1 _13096_ (.A(\cur_mb_mem[174][4] ),
    .B(_06046_),
    .C(_06758_),
    .X(_08141_));
 sky130_fd_sc_hd__and3_1 _13097_ (.A(\cur_mb_mem[187][4] ),
    .B(_06312_),
    .C(_06019_),
    .X(_08142_));
 sky130_fd_sc_hd__and3_1 _13098_ (.A(\cur_mb_mem[173][4] ),
    .B(_06762_),
    .C(_06755_),
    .X(_08143_));
 sky130_fd_sc_hd__a2111o_1 _13099_ (.A1(\cur_mb_mem[10][4] ),
    .A2(_06408_),
    .B1(_08141_),
    .C1(_08142_),
    .D1(_08143_),
    .X(_08144_));
 sky130_fd_sc_hd__and3_1 _13100_ (.A(\cur_mb_mem[233][4] ),
    .B(_06038_),
    .C(_06116_),
    .X(_08145_));
 sky130_fd_sc_hd__and3_1 _13101_ (.A(\cur_mb_mem[230][4] ),
    .B(_06204_),
    .C(_06255_),
    .X(_08146_));
 sky130_fd_sc_hd__and3_1 _13102_ (.A(\cur_mb_mem[63][4] ),
    .B(_06149_),
    .C(_06198_),
    .X(_08147_));
 sky130_fd_sc_hd__a2111o_2 _13103_ (.A1(\cur_mb_mem[231][4] ),
    .A2(_06180_),
    .B1(_08145_),
    .C1(_08146_),
    .D1(_08147_),
    .X(_08148_));
 sky130_fd_sc_hd__and3_1 _13104_ (.A(\cur_mb_mem[227][4] ),
    .B(_06289_),
    .C(_06766_),
    .X(_08149_));
 sky130_fd_sc_hd__and3_1 _13105_ (.A(\cur_mb_mem[224][4] ),
    .B(_06772_),
    .C(_06766_),
    .X(_08150_));
 sky130_fd_sc_hd__and3_1 _13106_ (.A(\cur_mb_mem[232][4] ),
    .B(_06832_),
    .C(_06918_),
    .X(_08151_));
 sky130_fd_sc_hd__a2111o_2 _13107_ (.A1(\cur_mb_mem[234][4] ),
    .A2(_06117_),
    .B1(_08149_),
    .C1(_08150_),
    .D1(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__or4_4 _13108_ (.A(_08140_),
    .B(_08144_),
    .C(_08148_),
    .D(_08152_),
    .X(_08153_));
 sky130_fd_sc_hd__or4_1 _13109_ (.A(_08102_),
    .B(_08119_),
    .C(_08136_),
    .D(_08153_),
    .X(_08154_));
 sky130_fd_sc_hd__and3_1 _13110_ (.A(\cur_mb_mem[154][4] ),
    .B(_06442_),
    .C(_06188_),
    .X(_08155_));
 sky130_fd_sc_hd__and3_1 _13111_ (.A(\cur_mb_mem[145][4] ),
    .B(_06188_),
    .C(_06076_),
    .X(_08156_));
 sky130_fd_sc_hd__and3_1 _13112_ (.A(\cur_mb_mem[100][4] ),
    .B(_06026_),
    .C(_06313_),
    .X(_08157_));
 sky130_fd_sc_hd__a2111o_1 _13113_ (.A1(\cur_mb_mem[159][4] ),
    .A2(_06174_),
    .B1(_08155_),
    .C1(_08156_),
    .D1(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__and3_1 _13114_ (.A(\cur_mb_mem[103][4] ),
    .B(_06267_),
    .C(_06851_),
    .X(_08159_));
 sky130_fd_sc_hd__and3_1 _13115_ (.A(\cur_mb_mem[99][4] ),
    .B(_06027_),
    .C(_06061_),
    .X(_08160_));
 sky130_fd_sc_hd__and3_1 _13116_ (.A(\cur_mb_mem[95][4] ),
    .B(_06120_),
    .C(_06378_),
    .X(_08161_));
 sky130_fd_sc_hd__a2111o_1 _13117_ (.A1(\cur_mb_mem[15][4] ),
    .A2(_06295_),
    .B1(_08159_),
    .C1(_08160_),
    .D1(_08161_),
    .X(_08162_));
 sky130_fd_sc_hd__and3_1 _13118_ (.A(\cur_mb_mem[105][4] ),
    .B(_05892_),
    .C(_06267_),
    .X(_08163_));
 sky130_fd_sc_hd__and3_1 _13119_ (.A(\cur_mb_mem[207][4] ),
    .B(_06099_),
    .C(_06789_),
    .X(_08164_));
 sky130_fd_sc_hd__and3_1 _13120_ (.A(\cur_mb_mem[96][4] ),
    .B(_06267_),
    .C(net236),
    .X(_08165_));
 sky130_fd_sc_hd__and3_1 _13121_ (.A(\cur_mb_mem[157][4] ),
    .B(_05944_),
    .C(_05977_),
    .X(_08166_));
 sky130_fd_sc_hd__or4_1 _13122_ (.A(_08163_),
    .B(_08164_),
    .C(_08165_),
    .D(_08166_),
    .X(_08167_));
 sky130_fd_sc_hd__and3_1 _13123_ (.A(\cur_mb_mem[101][4] ),
    .B(_05984_),
    .C(_06208_),
    .X(_08168_));
 sky130_fd_sc_hd__a221o_1 _13124_ (.A1(\cur_mb_mem[153][4] ),
    .A2(_06453_),
    .B1(_06305_),
    .B2(\cur_mb_mem[143][4] ),
    .C1(_08168_),
    .X(_08169_));
 sky130_fd_sc_hd__or4_2 _13125_ (.A(_08158_),
    .B(_08162_),
    .C(_08167_),
    .D(_08169_),
    .X(_08170_));
 sky130_fd_sc_hd__and3_1 _13126_ (.A(\cur_mb_mem[247][4] ),
    .B(_06032_),
    .C(_06851_),
    .X(_08171_));
 sky130_fd_sc_hd__and3_1 _13127_ (.A(\cur_mb_mem[202][4] ),
    .B(_06442_),
    .C(_06986_),
    .X(_08172_));
 sky130_fd_sc_hd__and3_1 _13128_ (.A(\cur_mb_mem[252][4] ),
    .B(_06158_),
    .C(_06422_),
    .X(_08173_));
 sky130_fd_sc_hd__a2111o_1 _13129_ (.A1(\cur_mb_mem[253][4] ),
    .A2(_06034_),
    .B1(_08171_),
    .C1(_08172_),
    .D1(_08173_),
    .X(_08174_));
 sky130_fd_sc_hd__and3_1 _13130_ (.A(\cur_mb_mem[212][4] ),
    .B(_06026_),
    .C(_06802_),
    .X(_08175_));
 sky130_fd_sc_hd__and3_1 _13131_ (.A(\cur_mb_mem[220][4] ),
    .B(_06321_),
    .C(_06802_),
    .X(_08176_));
 sky130_fd_sc_hd__and3_1 _13132_ (.A(\cur_mb_mem[104][4] ),
    .B(_06455_),
    .C(_06045_),
    .X(_08177_));
 sky130_fd_sc_hd__a2111o_1 _13133_ (.A1(\cur_mb_mem[250][4] ),
    .A2(_06443_),
    .B1(_08175_),
    .C1(_08176_),
    .D1(_08177_),
    .X(_08178_));
 sky130_fd_sc_hd__and3_1 _13134_ (.A(\cur_mb_mem[245][4] ),
    .B(_06032_),
    .C(_06131_),
    .X(_08179_));
 sky130_fd_sc_hd__and3_1 _13135_ (.A(\cur_mb_mem[193][4] ),
    .B(_06324_),
    .C(_05995_),
    .X(_08180_));
 sky130_fd_sc_hd__and3_4 _13136_ (.A(\cur_mb_mem[79][4] ),
    .B(_06120_),
    .C(_06233_),
    .X(_08181_));
 sky130_fd_sc_hd__a2111o_1 _13137_ (.A1(\cur_mb_mem[108][4] ),
    .A2(_06322_),
    .B1(_08179_),
    .C1(_08180_),
    .D1(_08181_),
    .X(_08182_));
 sky130_fd_sc_hd__and3_1 _13138_ (.A(\cur_mb_mem[197][4] ),
    .B(_06456_),
    .C(_06220_),
    .X(_08183_));
 sky130_fd_sc_hd__and3_1 _13139_ (.A(\cur_mb_mem[208][4] ),
    .B(_06270_),
    .C(_06009_),
    .X(_08184_));
 sky130_fd_sc_hd__and3_1 _13140_ (.A(\cur_mb_mem[205][4] ),
    .B(_06762_),
    .C(_06082_),
    .X(_08185_));
 sky130_fd_sc_hd__a2111o_1 _13141_ (.A1(\cur_mb_mem[111][4] ),
    .A2(_06069_),
    .B1(_08183_),
    .C1(_08184_),
    .D1(_08185_),
    .X(_08186_));
 sky130_fd_sc_hd__or4_4 _13142_ (.A(_08174_),
    .B(_08178_),
    .C(_08182_),
    .D(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__a32o_1 _13143_ (.A1(\cur_mb_mem[13][4] ),
    .A2(_06112_),
    .A3(_05946_),
    .B1(_06284_),
    .B2(\cur_mb_mem[162][4] ),
    .X(_08188_));
 sky130_fd_sc_hd__a32o_1 _13144_ (.A1(\cur_mb_mem[167][4] ),
    .A2(_06137_),
    .A3(_06097_),
    .B1(_06236_),
    .B2(\cur_mb_mem[21][4] ),
    .X(_08189_));
 sky130_fd_sc_hd__or2_1 _13145_ (.A(_08188_),
    .B(_08189_),
    .X(_08190_));
 sky130_fd_sc_hd__a32o_2 _13146_ (.A1(\cur_mb_mem[213][4] ),
    .A2(_05941_),
    .A3(_06132_),
    .B1(_06193_),
    .B2(\cur_mb_mem[166][4] ),
    .X(_08191_));
 sky130_fd_sc_hd__a32o_2 _13147_ (.A1(\cur_mb_mem[20][4] ),
    .A2(_05890_),
    .A3(_05975_),
    .B1(_06301_),
    .B2(\cur_mb_mem[11][4] ),
    .X(_08192_));
 sky130_fd_sc_hd__and3_1 _13148_ (.A(\cur_mb_mem[165][4] ),
    .B(_06825_),
    .C(_06220_),
    .X(_08193_));
 sky130_fd_sc_hd__and3_1 _13149_ (.A(\cur_mb_mem[6][4] ),
    .B(_06202_),
    .C(_06204_),
    .X(_08194_));
 sky130_fd_sc_hd__and3_1 _13150_ (.A(\cur_mb_mem[160][4] ),
    .B(_06192_),
    .C(_06772_),
    .X(_08195_));
 sky130_fd_sc_hd__a2111o_1 _13151_ (.A1(\cur_mb_mem[73][4] ),
    .A2(_06328_),
    .B1(_08193_),
    .C1(_08194_),
    .D1(_08195_),
    .X(_08196_));
 sky130_fd_sc_hd__and3_1 _13152_ (.A(\cur_mb_mem[186][4] ),
    .B(_05957_),
    .C(_06760_),
    .X(_08197_));
 sky130_fd_sc_hd__and3_1 _13153_ (.A(\cur_mb_mem[184][4] ),
    .B(_05982_),
    .C(_06830_),
    .X(_08198_));
 sky130_fd_sc_hd__and3_1 _13154_ (.A(\cur_mb_mem[185][4] ),
    .B(_06834_),
    .C(_06877_),
    .X(_08199_));
 sky130_fd_sc_hd__a2111o_1 _13155_ (.A1(\cur_mb_mem[74][4] ),
    .A2(_06417_),
    .B1(_08197_),
    .C1(_08198_),
    .D1(_08199_),
    .X(_08200_));
 sky130_fd_sc_hd__or4_1 _13156_ (.A(_08191_),
    .B(_08192_),
    .C(_08196_),
    .D(_08200_),
    .X(_08201_));
 sky130_fd_sc_hd__or4_1 _13157_ (.A(_08170_),
    .B(_08187_),
    .C(_08190_),
    .D(_08201_),
    .X(_08202_));
 sky130_fd_sc_hd__and3_1 _13158_ (.A(\cur_mb_mem[183][4] ),
    .B(_06013_),
    .C(_06851_),
    .X(_08203_));
 sky130_fd_sc_hd__and3_1 _13159_ (.A(\cur_mb_mem[131][4] ),
    .B(_06347_),
    .C(_05933_),
    .X(_08204_));
 sky130_fd_sc_hd__and3_1 _13160_ (.A(\cur_mb_mem[129][4] ),
    .B(_06353_),
    .C(_06382_),
    .X(_08205_));
 sky130_fd_sc_hd__a2111o_1 _13161_ (.A1(\cur_mb_mem[128][4] ),
    .A2(_06075_),
    .B1(_08203_),
    .C1(_08204_),
    .D1(_08205_),
    .X(_08206_));
 sky130_fd_sc_hd__and3_1 _13162_ (.A(\cur_mb_mem[182][4] ),
    .B(_06159_),
    .C(_06013_),
    .X(_08207_));
 sky130_fd_sc_hd__and3_1 _13163_ (.A(\cur_mb_mem[57][4] ),
    .B(_06849_),
    .C(_05909_),
    .X(_08208_));
 sky130_fd_sc_hd__and3_2 _13164_ (.A(\cur_mb_mem[107][4] ),
    .B(_06312_),
    .C(_06045_),
    .X(_08209_));
 sky130_fd_sc_hd__a2111o_1 _13165_ (.A1(\cur_mb_mem[135][4] ),
    .A2(_06462_),
    .B1(_08207_),
    .C1(_08208_),
    .D1(_08209_),
    .X(_08210_));
 sky130_fd_sc_hd__and3_1 _13166_ (.A(\cur_mb_mem[60][4] ),
    .B(_06849_),
    .C(_05901_),
    .X(_08211_));
 sky130_fd_sc_hd__and3_1 _13167_ (.A(\cur_mb_mem[55][4] ),
    .B(_06849_),
    .C(_06851_),
    .X(_08212_));
 sky130_fd_sc_hd__and3_1 _13168_ (.A(\cur_mb_mem[178][4] ),
    .B(_06079_),
    .C(_06018_),
    .X(_08213_));
 sky130_fd_sc_hd__and3_1 _13169_ (.A(\cur_mb_mem[177][4] ),
    .B(_06018_),
    .C(net230),
    .X(_08214_));
 sky130_fd_sc_hd__or4_1 _13170_ (.A(_08211_),
    .B(_08212_),
    .C(_08213_),
    .D(_08214_),
    .X(_08215_));
 sky130_fd_sc_hd__and3_1 _13171_ (.A(\cur_mb_mem[49][4] ),
    .B(_06350_),
    .C(_05995_),
    .X(_08216_));
 sky130_fd_sc_hd__and3_1 _13172_ (.A(\cur_mb_mem[36][4] ),
    .B(_06166_),
    .C(_06343_),
    .X(_08217_));
 sky130_fd_sc_hd__and3_1 _13173_ (.A(\cur_mb_mem[134][4] ),
    .B(_06199_),
    .C(_06146_),
    .X(_08218_));
 sky130_fd_sc_hd__a2111o_1 _13174_ (.A1(\cur_mb_mem[50][4] ),
    .A2(_06172_),
    .B1(_08216_),
    .C1(_08217_),
    .D1(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__or4_4 _13175_ (.A(_08206_),
    .B(_08210_),
    .C(_08215_),
    .D(_08219_),
    .X(_08220_));
 sky130_fd_sc_hd__and3_1 _13176_ (.A(\cur_mb_mem[31][4] ),
    .B(_06068_),
    .C(_06403_),
    .X(_08221_));
 sky130_fd_sc_hd__and3_2 _13177_ (.A(\cur_mb_mem[223][4] ),
    .B(_06068_),
    .C(_06348_),
    .X(_08222_));
 sky130_fd_sc_hd__and3_1 _13178_ (.A(\cur_mb_mem[163][4] ),
    .B(_06289_),
    .C(_06825_),
    .X(_08223_));
 sky130_fd_sc_hd__a2111o_1 _13179_ (.A1(\cur_mb_mem[47][4] ),
    .A2(_06259_),
    .B1(_08221_),
    .C1(_08222_),
    .D1(_08223_),
    .X(_08224_));
 sky130_fd_sc_hd__and3_2 _13180_ (.A(\cur_mb_mem[198][4] ),
    .B(_06159_),
    .C(_06986_),
    .X(_08225_));
 sky130_fd_sc_hd__and3_1 _13181_ (.A(\cur_mb_mem[102][4] ),
    .B(_06313_),
    .C(_06210_),
    .X(_08226_));
 sky130_fd_sc_hd__and3_1 _13182_ (.A(\cur_mb_mem[106][4] ),
    .B(_06115_),
    .C(_06045_),
    .X(_08227_));
 sky130_fd_sc_hd__a2111o_1 _13183_ (.A1(\cur_mb_mem[98][4] ),
    .A2(_06330_),
    .B1(_08225_),
    .C1(_08226_),
    .D1(_08227_),
    .X(_08228_));
 sky130_fd_sc_hd__and3_1 _13184_ (.A(\cur_mb_mem[175][4] ),
    .B(_06068_),
    .C(_06333_),
    .X(_08229_));
 sky130_fd_sc_hd__and3_1 _13185_ (.A(\cur_mb_mem[161][4] ),
    .B(_05995_),
    .C(_06758_),
    .X(_08230_));
 sky130_fd_sc_hd__and3_1 _13186_ (.A(\cur_mb_mem[180][4] ),
    .B(_06166_),
    .C(_06760_),
    .X(_08231_));
 sky130_fd_sc_hd__a2111o_1 _13187_ (.A1(\cur_mb_mem[97][4] ),
    .A2(_06077_),
    .B1(_08229_),
    .C1(_08230_),
    .D1(_08231_),
    .X(_08232_));
 sky130_fd_sc_hd__and3_1 _13188_ (.A(\cur_mb_mem[109][4] ),
    .B(_06045_),
    .C(_06490_),
    .X(_08233_));
 sky130_fd_sc_hd__and3_1 _13189_ (.A(\cur_mb_mem[148][4] ),
    .B(_06166_),
    .C(_06401_),
    .X(_08234_));
 sky130_fd_sc_hd__and3_1 _13190_ (.A(\cur_mb_mem[181][4] ),
    .B(_06830_),
    .C(_06794_),
    .X(_08235_));
 sky130_fd_sc_hd__a2111o_1 _13191_ (.A1(\cur_mb_mem[110][4] ),
    .A2(_06047_),
    .B1(_08233_),
    .C1(_08234_),
    .D1(_08235_),
    .X(_08236_));
 sky130_fd_sc_hd__or4_1 _13192_ (.A(_08224_),
    .B(_08228_),
    .C(_08232_),
    .D(_08236_),
    .X(_08237_));
 sky130_fd_sc_hd__and3_1 _13193_ (.A(\cur_mb_mem[48][4] ),
    .B(_06849_),
    .C(_06074_),
    .X(_08238_));
 sky130_fd_sc_hd__and3_1 _13194_ (.A(\cur_mb_mem[71][4] ),
    .B(_06143_),
    .C(_06461_),
    .X(_08239_));
 sky130_fd_sc_hd__and3_1 _13195_ (.A(\cur_mb_mem[64][4] ),
    .B(_06233_),
    .C(_06815_),
    .X(_08240_));
 sky130_fd_sc_hd__a2111o_1 _13196_ (.A1(\cur_mb_mem[65][4] ),
    .A2(_06483_),
    .B1(_08238_),
    .C1(_08239_),
    .D1(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__and3_1 _13197_ (.A(\cur_mb_mem[62][4] ),
    .B(_06849_),
    .C(_06366_),
    .X(_08242_));
 sky130_fd_sc_hd__and3_1 _13198_ (.A(\cur_mb_mem[58][4] ),
    .B(_06170_),
    .C(_05931_),
    .X(_08243_));
 sky130_fd_sc_hd__and3_1 _13199_ (.A(\cur_mb_mem[141][4] ),
    .B(_06490_),
    .C(_06842_),
    .X(_08244_));
 sky130_fd_sc_hd__a2111o_1 _13200_ (.A1(\cur_mb_mem[140][4] ),
    .A2(_06423_),
    .B1(_08242_),
    .C1(_08243_),
    .D1(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__and3_1 _13201_ (.A(\cur_mb_mem[44][4] ),
    .B(_06422_),
    .C(_06395_),
    .X(_08246_));
 sky130_fd_sc_hd__and3_1 _13202_ (.A(\cur_mb_mem[176][4] ),
    .B(_06039_),
    .C(_06009_),
    .X(_08247_));
 sky130_fd_sc_hd__and3_1 _13203_ (.A(\cur_mb_mem[56][4] ),
    .B(_06240_),
    .C(_06478_),
    .X(_08248_));
 sky130_fd_sc_hd__a2111o_2 _13204_ (.A1(\cur_mb_mem[61][4] ),
    .A2(_06359_),
    .B1(_08246_),
    .C1(_08247_),
    .D1(_08248_),
    .X(_08249_));
 sky130_fd_sc_hd__and3_1 _13205_ (.A(\cur_mb_mem[86][4] ),
    .B(_06931_),
    .C(_06140_),
    .X(_08250_));
 sky130_fd_sc_hd__and3_1 _13206_ (.A(\cur_mb_mem[93][4] ),
    .B(_05914_),
    .C(_06490_),
    .X(_08251_));
 sky130_fd_sc_hd__and3_1 _13207_ (.A(\cur_mb_mem[87][4] ),
    .B(_06927_),
    .C(_06896_),
    .X(_08252_));
 sky130_fd_sc_hd__a2111o_1 _13208_ (.A1(\cur_mb_mem[80][4] ),
    .A2(_06010_),
    .B1(_08250_),
    .C1(_08251_),
    .D1(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__or4_2 _13209_ (.A(_08241_),
    .B(_08245_),
    .C(_08249_),
    .D(_08253_),
    .X(_08254_));
 sky130_fd_sc_hd__and3_1 _13210_ (.A(\cur_mb_mem[235][4] ),
    .B(_06312_),
    .C(_06116_),
    .X(_08255_));
 sky130_fd_sc_hd__and3_1 _13211_ (.A(\cur_mb_mem[240][4] ),
    .B(_06165_),
    .C(_06815_),
    .X(_08256_));
 sky130_fd_sc_hd__and3_1 _13212_ (.A(\cur_mb_mem[249][4] ),
    .B(_06916_),
    .C(_06903_),
    .X(_08257_));
 sky130_fd_sc_hd__a2111o_1 _13213_ (.A1(\cur_mb_mem[248][4] ),
    .A2(_06411_),
    .B1(_08255_),
    .C1(_08256_),
    .D1(_08257_),
    .X(_08258_));
 sky130_fd_sc_hd__and3_1 _13214_ (.A(\cur_mb_mem[251][4] ),
    .B(_06158_),
    .C(_06312_),
    .X(_08259_));
 sky130_fd_sc_hd__and3_1 _13215_ (.A(\cur_mb_mem[59][4] ),
    .B(_06856_),
    .C(_06474_),
    .X(_08260_));
 sky130_fd_sc_hd__and3_1 _13216_ (.A(\cur_mb_mem[242][4] ),
    .B(_06916_),
    .C(_06080_),
    .X(_08261_));
 sky130_fd_sc_hd__a2111o_1 _13217_ (.A1(\cur_mb_mem[246][4] ),
    .A2(_06160_),
    .B1(_08259_),
    .C1(_08260_),
    .D1(_08261_),
    .X(_08262_));
 sky130_fd_sc_hd__and3_1 _13218_ (.A(\cur_mb_mem[228][4] ),
    .B(_06744_),
    .C(_06116_),
    .X(_08263_));
 sky130_fd_sc_hd__and3_1 _13219_ (.A(\cur_mb_mem[225][4] ),
    .B(_06841_),
    .C(_06766_),
    .X(_08264_));
 sky130_fd_sc_hd__and3_1 _13220_ (.A(\cur_mb_mem[254][4] ),
    .B(_06902_),
    .C(_06000_),
    .X(_08265_));
 sky130_fd_sc_hd__a2111o_1 _13221_ (.A1(\cur_mb_mem[255][4] ),
    .A2(_06304_),
    .B1(_08263_),
    .C1(_08264_),
    .D1(_08265_),
    .X(_08266_));
 sky130_fd_sc_hd__and3_1 _13222_ (.A(\cur_mb_mem[243][4] ),
    .B(_06916_),
    .C(_06770_),
    .X(_08267_));
 sky130_fd_sc_hd__and3_1 _13223_ (.A(\cur_mb_mem[226][4] ),
    .B(_06908_),
    .C(_06247_),
    .X(_08268_));
 sky130_fd_sc_hd__and3_1 _13224_ (.A(\cur_mb_mem[236][4] ),
    .B(_05902_),
    .C(_06775_),
    .X(_08269_));
 sky130_fd_sc_hd__a2111o_1 _13225_ (.A1(\cur_mb_mem[127][4] ),
    .A2(_06101_),
    .B1(_08267_),
    .C1(_08268_),
    .D1(_08269_),
    .X(_08270_));
 sky130_fd_sc_hd__or4_4 _13226_ (.A(_08258_),
    .B(_08262_),
    .C(_08266_),
    .D(_08270_),
    .X(_08271_));
 sky130_fd_sc_hd__or4_1 _13227_ (.A(_08220_),
    .B(_08237_),
    .C(_08254_),
    .D(_08271_),
    .X(_08272_));
 sky130_fd_sc_hd__and3_1 _13228_ (.A(\cur_mb_mem[94][4] ),
    .B(_06008_),
    .C(_06046_),
    .X(_08273_));
 sky130_fd_sc_hd__and3_1 _13229_ (.A(\cur_mb_mem[68][4] ),
    .B(_06744_),
    .C(_06121_),
    .X(_08274_));
 sky130_fd_sc_hd__and3_1 _13230_ (.A(\cur_mb_mem[91][4] ),
    .B(_06400_),
    .C(_05914_),
    .X(_08275_));
 sky130_fd_sc_hd__a2111o_1 _13231_ (.A1(\cur_mb_mem[136][4] ),
    .A2(_06292_),
    .B1(_08273_),
    .C1(_08274_),
    .D1(_08275_),
    .X(_08276_));
 sky130_fd_sc_hd__and3_1 _13232_ (.A(\cur_mb_mem[69][4] ),
    .B(_06143_),
    .C(_06220_),
    .X(_08277_));
 sky130_fd_sc_hd__and3_1 _13233_ (.A(\cur_mb_mem[90][4] ),
    .B(_06115_),
    .C(_06378_),
    .X(_08278_));
 sky130_fd_sc_hd__and3_4 _13234_ (.A(\cur_mb_mem[219][4] ),
    .B(_06400_),
    .C(_06814_),
    .X(_08279_));
 sky130_fd_sc_hd__a2111o_1 _13235_ (.A1(\cur_mb_mem[40][4] ),
    .A2(_06485_),
    .B1(_08277_),
    .C1(_08278_),
    .D1(_08279_),
    .X(_08280_));
 sky130_fd_sc_hd__and3_1 _13236_ (.A(\cur_mb_mem[46][4] ),
    .B(_06395_),
    .C(_06435_),
    .X(_08281_));
 sky130_fd_sc_hd__and3_1 _13237_ (.A(\cur_mb_mem[83][4] ),
    .B(_06931_),
    .C(_06289_),
    .X(_08282_));
 sky130_fd_sc_hd__and3_1 _13238_ (.A(\cur_mb_mem[92][4] ),
    .B(_06754_),
    .C(_06927_),
    .X(_08283_));
 sky130_fd_sc_hd__a2111o_1 _13239_ (.A1(\cur_mb_mem[70][4] ),
    .A2(_06144_),
    .B1(_08281_),
    .C1(_08282_),
    .D1(_08283_),
    .X(_08284_));
 sky130_fd_sc_hd__and3_1 _13240_ (.A(\cur_mb_mem[81][4] ),
    .B(_05914_),
    .C(_06841_),
    .X(_08285_));
 sky130_fd_sc_hd__and3_1 _13241_ (.A(\cur_mb_mem[82][4] ),
    .B(_06080_),
    .C(_06230_),
    .X(_08286_));
 sky130_fd_sc_hd__and3_1 _13242_ (.A(\cur_mb_mem[139][4] ),
    .B(_06942_),
    .C(_06859_),
    .X(_08287_));
 sky130_fd_sc_hd__a2111o_1 _13243_ (.A1(\cur_mb_mem[45][4] ),
    .A2(_06491_),
    .B1(_08285_),
    .C1(_08286_),
    .D1(_08287_),
    .X(_08288_));
 sky130_fd_sc_hd__or4_4 _13244_ (.A(_08276_),
    .B(_08280_),
    .C(_08284_),
    .D(_08288_),
    .X(_08289_));
 sky130_fd_sc_hd__and3_1 _13245_ (.A(\cur_mb_mem[130][4] ),
    .B(_06171_),
    .C(_06382_),
    .X(_08290_));
 sky130_fd_sc_hd__and3_1 _13246_ (.A(\cur_mb_mem[52][4] ),
    .B(_06350_),
    .C(_06744_),
    .X(_08291_));
 sky130_fd_sc_hd__and3_1 _13247_ (.A(\cur_mb_mem[54][4] ),
    .B(_06240_),
    .C(_06199_),
    .X(_08292_));
 sky130_fd_sc_hd__a2111o_4 _13248_ (.A1(\cur_mb_mem[53][4] ),
    .A2(_06221_),
    .B1(_08290_),
    .C1(_08291_),
    .D1(_08292_),
    .X(_08293_));
 sky130_fd_sc_hd__and3_1 _13249_ (.A(\cur_mb_mem[51][4] ),
    .B(_06170_),
    .C(_06355_),
    .X(_08294_));
 sky130_fd_sc_hd__and3_2 _13250_ (.A(\cur_mb_mem[229][4] ),
    .B(_06812_),
    .C(_06116_),
    .X(_08295_));
 sky130_fd_sc_hd__and3_1 _13251_ (.A(\cur_mb_mem[39][4] ),
    .B(_06343_),
    .C(_06708_),
    .X(_08296_));
 sky130_fd_sc_hd__a2111o_1 _13252_ (.A1(\cur_mb_mem[38][4] ),
    .A2(_06396_),
    .B1(_08294_),
    .C1(_08295_),
    .D1(_08296_),
    .X(_08297_));
 sky130_fd_sc_hd__and3_1 _13253_ (.A(\cur_mb_mem[191][4] ),
    .B(_06120_),
    .C(_06039_),
    .X(_08298_));
 sky130_fd_sc_hd__and3_1 _13254_ (.A(\cur_mb_mem[216][4] ),
    .B(_06455_),
    .C(_06814_),
    .X(_08299_));
 sky130_fd_sc_hd__and3_1 _13255_ (.A(\cur_mb_mem[37][4] ),
    .B(_06952_),
    .C(_06208_),
    .X(_08300_));
 sky130_fd_sc_hd__a2111o_1 _13256_ (.A1(\cur_mb_mem[239][4] ),
    .A2(_06125_),
    .B1(_08298_),
    .C1(_08299_),
    .D1(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__and3_2 _13257_ (.A(\cur_mb_mem[241][4] ),
    .B(_06165_),
    .C(_06841_),
    .X(_08302_));
 sky130_fd_sc_hd__and3_1 _13258_ (.A(\cur_mb_mem[218][4] ),
    .B(_06960_),
    .C(_06814_),
    .X(_08303_));
 sky130_fd_sc_hd__and3_1 _13259_ (.A(\cur_mb_mem[210][4] ),
    .B(_06380_),
    .C(_05947_),
    .X(_08304_));
 sky130_fd_sc_hd__a2111o_4 _13260_ (.A1(\cur_mb_mem[209][4] ),
    .A2(_06271_),
    .B1(_08302_),
    .C1(_08303_),
    .D1(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__or4_4 _13261_ (.A(_08293_),
    .B(_08297_),
    .C(_08301_),
    .D(_08305_),
    .X(_08306_));
 sky130_fd_sc_hd__and3_1 _13262_ (.A(\cur_mb_mem[214][4] ),
    .B(_06140_),
    .C(_06348_),
    .X(_08307_));
 sky130_fd_sc_hd__and3_1 _13263_ (.A(\cur_mb_mem[170][4] ),
    .B(_06115_),
    .C(_06825_),
    .X(_08308_));
 sky130_fd_sc_hd__and3_1 _13264_ (.A(\cur_mb_mem[199][4] ),
    .B(_06082_),
    .C(_06708_),
    .X(_08309_));
 sky130_fd_sc_hd__a2111o_2 _13265_ (.A1(\cur_mb_mem[200][4] ),
    .A2(_06457_),
    .B1(_08307_),
    .C1(_08308_),
    .D1(_08309_),
    .X(_08310_));
 sky130_fd_sc_hd__and3_1 _13266_ (.A(\cur_mb_mem[169][4] ),
    .B(_05892_),
    .C(_05921_),
    .X(_08311_));
 sky130_fd_sc_hd__and3_1 _13267_ (.A(\cur_mb_mem[222][4] ),
    .B(_05940_),
    .C(_05953_),
    .X(_08312_));
 sky130_fd_sc_hd__and3_1 _13268_ (.A(\cur_mb_mem[221][4] ),
    .B(_06033_),
    .C(_05940_),
    .X(_08313_));
 sky130_fd_sc_hd__and3_2 _13269_ (.A(\cur_mb_mem[32][4] ),
    .B(_06005_),
    .C(_06074_),
    .X(_08314_));
 sky130_fd_sc_hd__or4_4 _13270_ (.A(_08311_),
    .B(_08312_),
    .C(_08313_),
    .D(_08314_),
    .X(_08315_));
 sky130_fd_sc_hd__and3_1 _13271_ (.A(\cur_mb_mem[88][4] ),
    .B(_06455_),
    .C(_06931_),
    .X(_08316_));
 sky130_fd_sc_hd__and3_1 _13272_ (.A(\cur_mb_mem[137][4] ),
    .B(_06723_),
    .C(_06842_),
    .X(_08317_));
 sky130_fd_sc_hd__and3_1 _13273_ (.A(\cur_mb_mem[33][4] ),
    .B(_06087_),
    .C(_06912_),
    .X(_08318_));
 sky130_fd_sc_hd__a2111o_1 _13274_ (.A1(\cur_mb_mem[215][4] ),
    .A2(_06447_),
    .B1(_08316_),
    .C1(_08317_),
    .D1(_08318_),
    .X(_08319_));
 sky130_fd_sc_hd__and3_1 _13275_ (.A(\cur_mb_mem[89][4] ),
    .B(_06723_),
    .C(_06230_),
    .X(_08320_));
 sky130_fd_sc_hd__and3_1 _13276_ (.A(\cur_mb_mem[35][4] ),
    .B(_06980_),
    .C(_06952_),
    .X(_08321_));
 sky130_fd_sc_hd__and3_1 _13277_ (.A(\cur_mb_mem[138][4] ),
    .B(_05905_),
    .C(_06859_),
    .X(_08322_));
 sky130_fd_sc_hd__a2111o_1 _13278_ (.A1(\cur_mb_mem[34][4] ),
    .A2(_06393_),
    .B1(_08320_),
    .C1(_08321_),
    .D1(_08322_),
    .X(_08323_));
 sky130_fd_sc_hd__or4_1 _13279_ (.A(_08310_),
    .B(_08315_),
    .C(_08319_),
    .D(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__and3_2 _13280_ (.A(\cur_mb_mem[168][4] ),
    .B(net254),
    .C(_05921_),
    .X(_08325_));
 sky130_fd_sc_hd__and3_1 _13281_ (.A(\cur_mb_mem[194][4] ),
    .B(_06079_),
    .C(_06789_),
    .X(_08326_));
 sky130_fd_sc_hd__and3_1 _13282_ (.A(\cur_mb_mem[204][4] ),
    .B(_06321_),
    .C(_06986_),
    .X(_08327_));
 sky130_fd_sc_hd__and3_1 _13283_ (.A(\cur_mb_mem[211][4] ),
    .B(_06347_),
    .C(_06802_),
    .X(_08328_));
 sky130_fd_sc_hd__or4_1 _13284_ (.A(_08325_),
    .B(_08326_),
    .C(_08327_),
    .D(_08328_),
    .X(_08329_));
 sky130_fd_sc_hd__and3_1 _13285_ (.A(\cur_mb_mem[195][4] ),
    .B(_06061_),
    .C(_06789_),
    .X(_08330_));
 sky130_fd_sc_hd__and3_1 _13286_ (.A(\cur_mb_mem[142][4] ),
    .B(_05953_),
    .C(net244),
    .X(_08331_));
 sky130_fd_sc_hd__and3_1 _13287_ (.A(\cur_mb_mem[217][4] ),
    .B(_05909_),
    .C(_06802_),
    .X(_08332_));
 sky130_fd_sc_hd__and3_1 _13288_ (.A(\cur_mb_mem[201][4] ),
    .B(_05909_),
    .C(_06324_),
    .X(_08333_));
 sky130_fd_sc_hd__or4_1 _13289_ (.A(_08330_),
    .B(_08331_),
    .C(_08332_),
    .D(_08333_),
    .X(_08334_));
 sky130_fd_sc_hd__and3_1 _13290_ (.A(\cur_mb_mem[206][4] ),
    .B(_07075_),
    .C(_06082_),
    .X(_08335_));
 sky130_fd_sc_hd__and3_1 _13291_ (.A(\cur_mb_mem[192][4] ),
    .B(_06967_),
    .C(_06772_),
    .X(_08336_));
 sky130_fd_sc_hd__and3_2 _13292_ (.A(\cur_mb_mem[237][4] ),
    .B(_06246_),
    .C(_06775_),
    .X(_08337_));
 sky130_fd_sc_hd__a2111o_1 _13293_ (.A1(\cur_mb_mem[244][4] ),
    .A2(_06167_),
    .B1(_08335_),
    .C1(_08336_),
    .D1(_08337_),
    .X(_08338_));
 sky130_fd_sc_hd__and3_1 _13294_ (.A(\cur_mb_mem[171][4] ),
    .B(_06387_),
    .C(_07001_),
    .X(_08339_));
 sky130_fd_sc_hd__and3_1 _13295_ (.A(\cur_mb_mem[196][4] ),
    .B(_06215_),
    .C(_06997_),
    .X(_08340_));
 sky130_fd_sc_hd__and3_1 _13296_ (.A(\cur_mb_mem[238][4] ),
    .B(_07084_),
    .C(_06065_),
    .X(_08341_));
 sky130_fd_sc_hd__a2111o_1 _13297_ (.A1(\cur_mb_mem[203][4] ),
    .A2(_06325_),
    .B1(_08339_),
    .C1(_08340_),
    .D1(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__or4_4 _13298_ (.A(_08329_),
    .B(_08334_),
    .C(_08338_),
    .D(_08342_),
    .X(_08343_));
 sky130_fd_sc_hd__or4_1 _13299_ (.A(_08289_),
    .B(_08306_),
    .C(_08324_),
    .D(_08343_),
    .X(_08344_));
 sky130_fd_sc_hd__or4_4 _13300_ (.A(_08154_),
    .B(_08202_),
    .C(_08272_),
    .D(_08344_),
    .X(_08345_));
 sky130_fd_sc_hd__o22ai_4 _13301_ (.A1(\cur_mb_mem[0][4] ),
    .A2(_05908_),
    .B1(_08085_),
    .B2(_08345_),
    .Y(_08346_));
 sky130_fd_sc_hd__xor2_1 _13302_ (.A(net101),
    .B(_08346_),
    .X(_08347_));
 sky130_fd_sc_hd__and2_1 _13303_ (.A(_08074_),
    .B(_08347_),
    .X(_08348_));
 sky130_fd_sc_hd__a21boi_1 _13304_ (.A1(_08070_),
    .A2(_08073_),
    .B1_N(_08348_),
    .Y(_08349_));
 sky130_fd_sc_hd__nand2_1 _13305_ (.A(net102),
    .B(_07009_),
    .Y(_08350_));
 sky130_fd_sc_hd__nor2_1 _13306_ (.A(net101),
    .B(_08346_),
    .Y(_08351_));
 sky130_fd_sc_hd__and2_1 _13307_ (.A(_08350_),
    .B(_08351_),
    .X(_08352_));
 sky130_fd_sc_hd__or2_1 _13308_ (.A(\cur_mb_mem[0][6] ),
    .B(_05908_),
    .X(_08353_));
 sky130_fd_sc_hd__or2_1 _13309_ (.A(_06514_),
    .B(_06679_),
    .X(_08354_));
 sky130_fd_sc_hd__a21o_1 _13310_ (.A1(_08353_),
    .A2(_08354_),
    .B1(_06680_),
    .X(_08355_));
 sky130_fd_sc_hd__o41a_2 _13311_ (.A1(_06681_),
    .A2(_07010_),
    .A3(_08349_),
    .A4(_08352_),
    .B1(_08355_),
    .X(_08356_));
 sky130_fd_sc_hd__and2_1 _13312_ (.A(_06498_),
    .B(_08356_),
    .X(_08357_));
 sky130_fd_sc_hd__inv_2 _13313_ (.A(_08355_),
    .Y(_08358_));
 sky130_fd_sc_hd__and2_1 _13314_ (.A(net98),
    .B(_07286_),
    .X(_08359_));
 sky130_fd_sc_hd__nor2_1 _13315_ (.A(net98),
    .B(_07286_),
    .Y(_08360_));
 sky130_fd_sc_hd__nor2_1 _13316_ (.A(net97),
    .B(_07551_),
    .Y(_08361_));
 sky130_fd_sc_hd__nor2_1 _13317_ (.A(_08360_),
    .B(_08361_),
    .Y(_08362_));
 sky130_fd_sc_hd__nor2_1 _13318_ (.A(_08359_),
    .B(_08362_),
    .Y(_08363_));
 sky130_fd_sc_hd__o21ai_1 _13319_ (.A1(_07820_),
    .A2(net211),
    .B1(net99),
    .Y(_08364_));
 sky130_fd_sc_hd__o21a_1 _13320_ (.A1(_08068_),
    .A2(_08363_),
    .B1(_08364_),
    .X(_08365_));
 sky130_fd_sc_hd__o21a_1 _13321_ (.A1(_08072_),
    .A2(_08365_),
    .B1(_08071_),
    .X(_08366_));
 sky130_fd_sc_hd__nand2_1 _13322_ (.A(net101),
    .B(_08346_),
    .Y(_08367_));
 sky130_fd_sc_hd__o21a_1 _13323_ (.A1(_08351_),
    .A2(_08366_),
    .B1(_08367_),
    .X(_08368_));
 sky130_fd_sc_hd__o21a_1 _13324_ (.A1(_07010_),
    .A2(_08368_),
    .B1(_08350_),
    .X(_08369_));
 sky130_fd_sc_hd__nor2_1 _13325_ (.A(_06681_),
    .B(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__nor2_1 _13326_ (.A(_08068_),
    .B(_08069_),
    .Y(_08371_));
 sky130_fd_sc_hd__and2b_1 _13327_ (.A_N(_07819_),
    .B(_08371_),
    .X(_08372_));
 sky130_fd_sc_hd__and4bb_1 _13328_ (.A_N(_07552_),
    .B_N(_06681_),
    .C(_08348_),
    .D(_08362_),
    .X(_08373_));
 sky130_fd_sc_hd__and2_1 _13329_ (.A(net104),
    .B(_06497_),
    .X(_08374_));
 sky130_fd_sc_hd__a21oi_2 _13330_ (.A1(_08372_),
    .A2(_08373_),
    .B1(_08374_),
    .Y(_08375_));
 sky130_fd_sc_hd__a21o_1 _13331_ (.A1(_08356_),
    .A2(_08375_),
    .B1(_06498_),
    .X(_08376_));
 sky130_fd_sc_hd__o31a_1 _13332_ (.A1(_08358_),
    .A2(_08370_),
    .A3(_08376_),
    .B1(_08374_),
    .X(_08377_));
 sky130_fd_sc_hd__o21a_1 _13333_ (.A1(_08357_),
    .A2(_08377_),
    .B1(\current_accum_sad[7] ),
    .X(_08378_));
 sky130_fd_sc_hd__nor3_1 _13334_ (.A(\current_accum_sad[7] ),
    .B(_08357_),
    .C(_08377_),
    .Y(_08379_));
 sky130_fd_sc_hd__nor2_1 _13335_ (.A(_08378_),
    .B(_08379_),
    .Y(_08380_));
 sky130_fd_sc_hd__nand2_1 _13336_ (.A(_08070_),
    .B(_08073_),
    .Y(_08381_));
 sky130_fd_sc_hd__a21oi_1 _13337_ (.A1(_08367_),
    .A2(_08381_),
    .B1(_08351_),
    .Y(_08382_));
 sky130_fd_sc_hd__mux2_1 _13338_ (.A0(_08368_),
    .A1(_08382_),
    .S(_08376_),
    .X(_08383_));
 sky130_fd_sc_hd__xnor2_1 _13339_ (.A(_08074_),
    .B(_08383_),
    .Y(_08384_));
 sky130_fd_sc_hd__or2_1 _13340_ (.A(\current_accum_sad[5] ),
    .B(_08384_),
    .X(_08385_));
 sky130_fd_sc_hd__a21oi_4 _13341_ (.A1(_08356_),
    .A2(_08375_),
    .B1(_06498_),
    .Y(_08386_));
 sky130_fd_sc_hd__nand2_1 _13342_ (.A(_08366_),
    .B(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__o21ai_1 _13343_ (.A1(_08381_),
    .A2(_08386_),
    .B1(_08387_),
    .Y(_08388_));
 sky130_fd_sc_hd__xnor2_1 _13344_ (.A(_08347_),
    .B(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__or2_1 _13345_ (.A(\current_accum_sad[4] ),
    .B(_08389_),
    .X(_08390_));
 sky130_fd_sc_hd__nand2_1 _13346_ (.A(_07552_),
    .B(_07553_),
    .Y(_08391_));
 sky130_fd_sc_hd__o21ai_1 _13347_ (.A1(_08068_),
    .A2(_08391_),
    .B1(_08364_),
    .Y(_08392_));
 sky130_fd_sc_hd__mux2_1 _13348_ (.A0(_08365_),
    .A1(_08392_),
    .S(_08376_),
    .X(_08393_));
 sky130_fd_sc_hd__xor2_1 _13349_ (.A(_07819_),
    .B(_08393_),
    .X(_08394_));
 sky130_fd_sc_hd__or2_1 _13350_ (.A(\current_accum_sad[3] ),
    .B(_08394_),
    .X(_08395_));
 sky130_fd_sc_hd__inv_2 _13351_ (.A(_08391_),
    .Y(_08396_));
 sky130_fd_sc_hd__mux2_1 _13352_ (.A0(_08396_),
    .A1(_08363_),
    .S(_08386_),
    .X(_08397_));
 sky130_fd_sc_hd__xnor2_1 _13353_ (.A(_08371_),
    .B(_08397_),
    .Y(_08398_));
 sky130_fd_sc_hd__xor2_1 _13354_ (.A(\current_accum_sad[2] ),
    .B(_08398_),
    .X(_08399_));
 sky130_fd_sc_hd__and2_1 _13355_ (.A(net97),
    .B(_07551_),
    .X(_08400_));
 sky130_fd_sc_hd__o21a_1 _13356_ (.A1(_08400_),
    .A2(_08361_),
    .B1(\current_accum_sad[0] ),
    .X(_08401_));
 sky130_fd_sc_hd__inv_2 _13357_ (.A(_08401_),
    .Y(_08402_));
 sky130_fd_sc_hd__inv_2 _13358_ (.A(\current_accum_sad[1] ),
    .Y(_08403_));
 sky130_fd_sc_hd__nor2_1 _13359_ (.A(_08359_),
    .B(_08360_),
    .Y(_08404_));
 sky130_fd_sc_hd__a211o_1 _13360_ (.A1(_08356_),
    .A2(_08375_),
    .B1(_08361_),
    .C1(_06498_),
    .X(_08405_));
 sky130_fd_sc_hd__o211ai_1 _13361_ (.A1(_08400_),
    .A2(_08386_),
    .B1(_08404_),
    .C1(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__a2111oi_1 _13362_ (.A1(_08356_),
    .A2(_08375_),
    .B1(net97),
    .C1(_06498_),
    .D1(_07551_),
    .Y(_08407_));
 sky130_fd_sc_hd__a211o_1 _13363_ (.A1(_08400_),
    .A2(_08376_),
    .B1(_08404_),
    .C1(_08407_),
    .X(_08408_));
 sky130_fd_sc_hd__and3_1 _13364_ (.A(_08403_),
    .B(_08406_),
    .C(_08408_),
    .X(_08409_));
 sky130_fd_sc_hd__a21oi_1 _13365_ (.A1(_08406_),
    .A2(_08408_),
    .B1(_08403_),
    .Y(_08410_));
 sky130_fd_sc_hd__o21bai_2 _13366_ (.A1(_08402_),
    .A2(_08409_),
    .B1_N(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__and2_1 _13367_ (.A(\current_accum_sad[2] ),
    .B(_08398_),
    .X(_08412_));
 sky130_fd_sc_hd__a21o_1 _13368_ (.A1(_08399_),
    .A2(_08411_),
    .B1(_08412_),
    .X(_08413_));
 sky130_fd_sc_hd__and2_1 _13369_ (.A(\current_accum_sad[3] ),
    .B(_08394_),
    .X(_08414_));
 sky130_fd_sc_hd__a21o_1 _13370_ (.A1(_08395_),
    .A2(_08413_),
    .B1(_08414_),
    .X(_08415_));
 sky130_fd_sc_hd__and2_1 _13371_ (.A(\current_accum_sad[4] ),
    .B(_08389_),
    .X(_08416_));
 sky130_fd_sc_hd__a21o_1 _13372_ (.A1(_08390_),
    .A2(_08415_),
    .B1(_08416_),
    .X(_08417_));
 sky130_fd_sc_hd__and2_1 _13373_ (.A(\current_accum_sad[5] ),
    .B(_08384_),
    .X(_08418_));
 sky130_fd_sc_hd__a21o_1 _13374_ (.A1(_08385_),
    .A2(_08417_),
    .B1(_08418_),
    .X(_08419_));
 sky130_fd_sc_hd__inv_2 _13375_ (.A(\current_accum_sad[6] ),
    .Y(_08420_));
 sky130_fd_sc_hd__nor2_1 _13376_ (.A(_08358_),
    .B(_06681_),
    .Y(_08421_));
 sky130_fd_sc_hd__nand2_1 _13377_ (.A(_08369_),
    .B(_08386_),
    .Y(_08422_));
 sky130_fd_sc_hd__o41a_1 _13378_ (.A1(_07010_),
    .A2(_08349_),
    .A3(_08352_),
    .A4(_08386_),
    .B1(_08422_),
    .X(_08423_));
 sky130_fd_sc_hd__xnor2_1 _13379_ (.A(_08421_),
    .B(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__nor2_1 _13380_ (.A(_08420_),
    .B(_08424_),
    .Y(_08425_));
 sky130_fd_sc_hd__and2_1 _13381_ (.A(_08420_),
    .B(_08424_),
    .X(_08426_));
 sky130_fd_sc_hd__nor2_1 _13382_ (.A(_08425_),
    .B(_08426_),
    .Y(_08427_));
 sky130_fd_sc_hd__a21o_1 _13383_ (.A1(_08419_),
    .A2(_08427_),
    .B1(_08425_),
    .X(_08428_));
 sky130_fd_sc_hd__a21o_1 _13384_ (.A1(_08380_),
    .A2(_08428_),
    .B1(_08378_),
    .X(_08429_));
 sky130_fd_sc_hd__and4_1 _13385_ (.A(\current_accum_sad[10] ),
    .B(\current_accum_sad[9] ),
    .C(\current_accum_sad[8] ),
    .D(_08429_),
    .X(_08430_));
 sky130_fd_sc_hd__and3_1 _13386_ (.A(\current_accum_sad[12] ),
    .B(\current_accum_sad[11] ),
    .C(_08430_),
    .X(_08431_));
 sky130_fd_sc_hd__and2_1 _13387_ (.A(\current_accum_sad[13] ),
    .B(_08431_),
    .X(_08432_));
 sky130_fd_sc_hd__nand2_1 _13388_ (.A(\current_accum_sad[14] ),
    .B(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__xor2_1 _13389_ (.A(\current_accum_sad[15] ),
    .B(_08433_),
    .X(_08434_));
 sky130_fd_sc_hd__and2_1 _13390_ (.A(_05886_),
    .B(_08434_),
    .X(_08435_));
 sky130_fd_sc_hd__or2_1 _13391_ (.A(\current_accum_sad[14] ),
    .B(_08432_),
    .X(_08436_));
 sky130_fd_sc_hd__inv_2 _13392_ (.A(net217),
    .Y(_08437_));
 sky130_fd_sc_hd__a21oi_2 _13393_ (.A1(_08433_),
    .A2(_08436_),
    .B1(_08437_),
    .Y(_08438_));
 sky130_fd_sc_hd__nor2_1 _13394_ (.A(\current_accum_sad[13] ),
    .B(_08431_),
    .Y(_08439_));
 sky130_fd_sc_hd__or2_1 _13395_ (.A(_08432_),
    .B(_08439_),
    .X(_08440_));
 sky130_fd_sc_hd__and2_1 _13396_ (.A(_05886_),
    .B(_08440_),
    .X(_08441_));
 sky130_fd_sc_hd__a21oi_1 _13397_ (.A1(\current_accum_sad[11] ),
    .A2(_08430_),
    .B1(\current_accum_sad[12] ),
    .Y(_08442_));
 sky130_fd_sc_hd__or2_1 _13398_ (.A(_08431_),
    .B(_08442_),
    .X(_08443_));
 sky130_fd_sc_hd__and2_1 _13399_ (.A(_05886_),
    .B(_08443_),
    .X(_08444_));
 sky130_fd_sc_hd__inv_2 _13400_ (.A(\min_sad_reg[11] ),
    .Y(_08445_));
 sky130_fd_sc_hd__xnor2_1 _13401_ (.A(\current_accum_sad[11] ),
    .B(_08430_),
    .Y(_08446_));
 sky130_fd_sc_hd__nand2_1 _13402_ (.A(_05886_),
    .B(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__a2bb2o_1 _13403_ (.A1_N(_08445_),
    .A2_N(_08447_),
    .B1(_08444_),
    .B2(\min_sad_reg[12] ),
    .X(_08448_));
 sky130_fd_sc_hd__inv_2 _13404_ (.A(\min_sad_reg[9] ),
    .Y(_08449_));
 sky130_fd_sc_hd__nand3_1 _13405_ (.A(\current_accum_sad[9] ),
    .B(\current_accum_sad[8] ),
    .C(_08429_),
    .Y(_08450_));
 sky130_fd_sc_hd__a21o_1 _13406_ (.A1(\current_accum_sad[8] ),
    .A2(_08429_),
    .B1(\current_accum_sad[9] ),
    .X(_08451_));
 sky130_fd_sc_hd__a21o_1 _13407_ (.A1(_08450_),
    .A2(_08451_),
    .B1(_08437_),
    .X(_08452_));
 sky130_fd_sc_hd__inv_2 _13408_ (.A(\min_sad_reg[8] ),
    .Y(_08453_));
 sky130_fd_sc_hd__nand2_1 _13409_ (.A(\current_accum_sad[8] ),
    .B(_08429_),
    .Y(_08454_));
 sky130_fd_sc_hd__or2_1 _13410_ (.A(\current_accum_sad[8] ),
    .B(_08429_),
    .X(_08455_));
 sky130_fd_sc_hd__a21o_1 _13411_ (.A1(_08454_),
    .A2(_08455_),
    .B1(_08437_),
    .X(_08456_));
 sky130_fd_sc_hd__or2_1 _13412_ (.A(_08453_),
    .B(_08456_),
    .X(_08457_));
 sky130_fd_sc_hd__inv_2 _13413_ (.A(\min_sad_reg[7] ),
    .Y(_08458_));
 sky130_fd_sc_hd__nand2_1 _13414_ (.A(_08380_),
    .B(_08428_),
    .Y(_08459_));
 sky130_fd_sc_hd__or2_1 _13415_ (.A(_08380_),
    .B(_08428_),
    .X(_08460_));
 sky130_fd_sc_hd__a21o_1 _13416_ (.A1(_08459_),
    .A2(_08460_),
    .B1(_08437_),
    .X(_08461_));
 sky130_fd_sc_hd__xnor2_1 _13417_ (.A(_08419_),
    .B(_08427_),
    .Y(_08462_));
 sky130_fd_sc_hd__nand2_1 _13418_ (.A(net217),
    .B(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__inv_2 _13419_ (.A(\min_sad_reg[6] ),
    .Y(_08464_));
 sky130_fd_sc_hd__or2b_1 _13420_ (.A(_08418_),
    .B_N(_08385_),
    .X(_08465_));
 sky130_fd_sc_hd__xor2_2 _13421_ (.A(_08465_),
    .B(_08417_),
    .X(_08466_));
 sky130_fd_sc_hd__a21o_1 _13422_ (.A1(net217),
    .A2(_08466_),
    .B1(\min_sad_reg[5] ),
    .X(_08467_));
 sky130_fd_sc_hd__inv_2 _13423_ (.A(\min_sad_reg[4] ),
    .Y(_08468_));
 sky130_fd_sc_hd__or2b_1 _13424_ (.A(_08416_),
    .B_N(_08390_),
    .X(_08469_));
 sky130_fd_sc_hd__xor2_1 _13425_ (.A(_08469_),
    .B(_08415_),
    .X(_08470_));
 sky130_fd_sc_hd__nand2_1 _13426_ (.A(net217),
    .B(_08470_),
    .Y(_08471_));
 sky130_fd_sc_hd__nand2_1 _13427_ (.A(_08468_),
    .B(_08471_),
    .Y(_08472_));
 sky130_fd_sc_hd__inv_2 _13428_ (.A(\min_sad_reg[2] ),
    .Y(_08473_));
 sky130_fd_sc_hd__xnor2_1 _13429_ (.A(_08399_),
    .B(_08411_),
    .Y(_08474_));
 sky130_fd_sc_hd__nand2_2 _13430_ (.A(net217),
    .B(_08474_),
    .Y(_08475_));
 sky130_fd_sc_hd__or2_1 _13431_ (.A(_08410_),
    .B(_08409_),
    .X(_08476_));
 sky130_fd_sc_hd__xnor2_1 _13432_ (.A(_08402_),
    .B(_08476_),
    .Y(_08477_));
 sky130_fd_sc_hd__nand2_1 _13433_ (.A(net217),
    .B(_08477_),
    .Y(_08478_));
 sky130_fd_sc_hd__or3_1 _13434_ (.A(\current_accum_sad[0] ),
    .B(_08400_),
    .C(_08361_),
    .X(_08479_));
 sky130_fd_sc_hd__and2_1 _13435_ (.A(_08402_),
    .B(_08479_),
    .X(_08480_));
 sky130_fd_sc_hd__and3b_1 _13436_ (.A_N(_08480_),
    .B(net217),
    .C(\min_sad_reg[0] ),
    .X(_08481_));
 sky130_fd_sc_hd__nor2_1 _13437_ (.A(\min_sad_reg[1] ),
    .B(_08481_),
    .Y(_08482_));
 sky130_fd_sc_hd__nand2_1 _13438_ (.A(\min_sad_reg[1] ),
    .B(_08481_),
    .Y(_08483_));
 sky130_fd_sc_hd__o221a_1 _13439_ (.A1(_08473_),
    .A2(_08475_),
    .B1(_08478_),
    .B2(_08482_),
    .C1(_08483_),
    .X(_08484_));
 sky130_fd_sc_hd__inv_2 _13440_ (.A(\min_sad_reg[3] ),
    .Y(_08485_));
 sky130_fd_sc_hd__or2b_1 _13441_ (.A(_08414_),
    .B_N(_08395_),
    .X(_08486_));
 sky130_fd_sc_hd__xor2_1 _13442_ (.A(_08486_),
    .B(_08413_),
    .X(_08487_));
 sky130_fd_sc_hd__nand2_1 _13443_ (.A(net217),
    .B(_08487_),
    .Y(_08488_));
 sky130_fd_sc_hd__a22o_1 _13444_ (.A1(_08485_),
    .A2(_08488_),
    .B1(_08475_),
    .B2(_08473_),
    .X(_08489_));
 sky130_fd_sc_hd__or2_1 _13445_ (.A(_08485_),
    .B(_08488_),
    .X(_08490_));
 sky130_fd_sc_hd__o221ai_1 _13446_ (.A1(_08468_),
    .A2(_08471_),
    .B1(_08484_),
    .B2(_08489_),
    .C1(_08490_),
    .Y(_08491_));
 sky130_fd_sc_hd__a32o_1 _13447_ (.A1(\min_sad_reg[5] ),
    .A2(net217),
    .A3(_08466_),
    .B1(_08472_),
    .B2(_08491_),
    .X(_08492_));
 sky130_fd_sc_hd__o2bb2a_1 _13448_ (.A1_N(_08467_),
    .A2_N(_08492_),
    .B1(_08464_),
    .B2(_08463_),
    .X(_08493_));
 sky130_fd_sc_hd__a221o_1 _13449_ (.A1(_08458_),
    .A2(_08461_),
    .B1(_08463_),
    .B2(_08464_),
    .C1(_08493_),
    .X(_08494_));
 sky130_fd_sc_hd__o21a_1 _13450_ (.A1(_08458_),
    .A2(_08461_),
    .B1(_08494_),
    .X(_08495_));
 sky130_fd_sc_hd__and2_1 _13451_ (.A(_08453_),
    .B(_08456_),
    .X(_08496_));
 sky130_fd_sc_hd__a221o_1 _13452_ (.A1(_08449_),
    .A2(_08452_),
    .B1(_08457_),
    .B2(_08495_),
    .C1(_08496_),
    .X(_08497_));
 sky130_fd_sc_hd__a21oi_1 _13453_ (.A1(_08450_),
    .A2(_08451_),
    .B1(_08437_),
    .Y(_08498_));
 sky130_fd_sc_hd__xor2_1 _13454_ (.A(\current_accum_sad[10] ),
    .B(_08450_),
    .X(_08499_));
 sky130_fd_sc_hd__and2_1 _13455_ (.A(_05886_),
    .B(_08499_),
    .X(_08500_));
 sky130_fd_sc_hd__a22oi_1 _13456_ (.A1(\min_sad_reg[9] ),
    .A2(_08498_),
    .B1(_08500_),
    .B2(\min_sad_reg[10] ),
    .Y(_08501_));
 sky130_fd_sc_hd__a2bb2o_1 _13457_ (.A1_N(\min_sad_reg[10] ),
    .A2_N(_08500_),
    .B1(_08447_),
    .B2(_08445_),
    .X(_08502_));
 sky130_fd_sc_hd__a21oi_1 _13458_ (.A1(_08497_),
    .A2(_08501_),
    .B1(_08502_),
    .Y(_08503_));
 sky130_fd_sc_hd__o22a_1 _13459_ (.A1(\min_sad_reg[12] ),
    .A2(_08444_),
    .B1(_08448_),
    .B2(_08503_),
    .X(_08504_));
 sky130_fd_sc_hd__a221o_1 _13460_ (.A1(\min_sad_reg[14] ),
    .A2(_08438_),
    .B1(_08441_),
    .B2(\min_sad_reg[13] ),
    .C1(_08504_),
    .X(_08505_));
 sky130_fd_sc_hd__a211o_1 _13461_ (.A1(\min_sad_reg[14] ),
    .A2(_08438_),
    .B1(_08441_),
    .C1(\min_sad_reg[13] ),
    .X(_08506_));
 sky130_fd_sc_hd__o221a_1 _13462_ (.A1(\min_sad_reg[15] ),
    .A2(_08435_),
    .B1(_08438_),
    .B2(\min_sad_reg[14] ),
    .C1(_08506_),
    .X(_08507_));
 sky130_fd_sc_hd__a22oi_4 _13463_ (.A1(\min_sad_reg[15] ),
    .A2(_08435_),
    .B1(_08505_),
    .B2(_08507_),
    .Y(_08508_));
 sky130_fd_sc_hd__a21o_1 _13464_ (.A1(\state[3] ),
    .A2(shex_load),
    .B1(_04442_),
    .X(_08509_));
 sky130_fd_sc_hd__or4b_4 _13465_ (.A(_04686_),
    .B(_08508_),
    .C(_08509_),
    .D_N(net266),
    .X(_08510_));
 sky130_fd_sc_hd__buf_4 _13466_ (.A(_08510_),
    .X(_08511_));
 sky130_fd_sc_hd__mux2_1 _13467_ (.A0(\cand_x[0] ),
    .A1(\best_cand_x[0] ),
    .S(_08511_),
    .X(_08512_));
 sky130_fd_sc_hd__clkbuf_1 _13468_ (.A(_08512_),
    .X(_00008_));
 sky130_fd_sc_hd__mux2_1 _13469_ (.A0(\cand_x[1] ),
    .A1(net1597),
    .S(_08511_),
    .X(_08513_));
 sky130_fd_sc_hd__clkbuf_1 _13470_ (.A(_08513_),
    .X(_00009_));
 sky130_fd_sc_hd__mux2_1 _13471_ (.A0(\cand_x[2] ),
    .A1(net1839),
    .S(_08511_),
    .X(_08514_));
 sky130_fd_sc_hd__clkbuf_1 _13472_ (.A(_08514_),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _13473_ (.A0(net1996),
    .A1(net1602),
    .S(_08511_),
    .X(_08515_));
 sky130_fd_sc_hd__clkbuf_1 _13474_ (.A(_08515_),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _13475_ (.A0(\cand_x[4] ),
    .A1(net1787),
    .S(_08511_),
    .X(_08516_));
 sky130_fd_sc_hd__clkbuf_1 _13476_ (.A(_08516_),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _13477_ (.A0(\cand_x[5] ),
    .A1(net1845),
    .S(_08511_),
    .X(_08517_));
 sky130_fd_sc_hd__clkbuf_1 _13478_ (.A(_08517_),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _13479_ (.A0(_04475_),
    .A1(net565),
    .S(_08511_),
    .X(_08518_));
 sky130_fd_sc_hd__clkbuf_1 _13480_ (.A(_08518_),
    .X(_00014_));
 sky130_fd_sc_hd__or2_1 _13481_ (.A(_08437_),
    .B(_08480_),
    .X(_08519_));
 sky130_fd_sc_hd__a21o_4 _13482_ (.A1(_04463_),
    .A2(_08508_),
    .B1(_08509_),
    .X(_08520_));
 sky130_fd_sc_hd__clkbuf_4 _13483_ (.A(_08520_),
    .X(_08521_));
 sky130_fd_sc_hd__a21oi_4 _13484_ (.A1(_04956_),
    .A2(_04686_),
    .B1(_08520_),
    .Y(_08522_));
 sky130_fd_sc_hd__clkbuf_4 _13485_ (.A(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__o32a_1 _13486_ (.A1(_04689_),
    .A2(_08519_),
    .A3(_08521_),
    .B1(_08523_),
    .B2(net1934),
    .X(_00015_));
 sky130_fd_sc_hd__o32a_1 _13487_ (.A1(_04689_),
    .A2(_08478_),
    .A3(_08521_),
    .B1(_08523_),
    .B2(net1973),
    .X(_00016_));
 sky130_fd_sc_hd__o32a_1 _13488_ (.A1(_04689_),
    .A2(_08475_),
    .A3(_08521_),
    .B1(_08523_),
    .B2(net1767),
    .X(_00017_));
 sky130_fd_sc_hd__o32a_1 _13489_ (.A1(_04689_),
    .A2(_08488_),
    .A3(_08521_),
    .B1(_08523_),
    .B2(net1511),
    .X(_00018_));
 sky130_fd_sc_hd__o32a_1 _13490_ (.A1(_04689_),
    .A2(_08471_),
    .A3(_08521_),
    .B1(_08523_),
    .B2(net1459),
    .X(_00019_));
 sky130_fd_sc_hd__nand2_1 _13491_ (.A(_05886_),
    .B(_08466_),
    .Y(_08524_));
 sky130_fd_sc_hd__o32a_1 _13492_ (.A1(_04689_),
    .A2(_08524_),
    .A3(_08521_),
    .B1(_08523_),
    .B2(net1774),
    .X(_00020_));
 sky130_fd_sc_hd__o32a_1 _13493_ (.A1(_04689_),
    .A2(_08463_),
    .A3(_08521_),
    .B1(_08523_),
    .B2(net1599),
    .X(_00021_));
 sky130_fd_sc_hd__o32a_1 _13494_ (.A1(_04689_),
    .A2(_08461_),
    .A3(_08521_),
    .B1(_08523_),
    .B2(\min_sad_reg[7] ),
    .X(_00022_));
 sky130_fd_sc_hd__o32a_1 _13495_ (.A1(_04689_),
    .A2(_08456_),
    .A3(_08521_),
    .B1(_08523_),
    .B2(net1402),
    .X(_00023_));
 sky130_fd_sc_hd__o32a_1 _13496_ (.A1(_05485_),
    .A2(_08452_),
    .A3(_08521_),
    .B1(_08523_),
    .B2(net1832),
    .X(_00024_));
 sky130_fd_sc_hd__nand2_1 _13497_ (.A(_05886_),
    .B(_08499_),
    .Y(_08525_));
 sky130_fd_sc_hd__o32a_1 _13498_ (.A1(_05485_),
    .A2(_08525_),
    .A3(_08520_),
    .B1(_08522_),
    .B2(\min_sad_reg[10] ),
    .X(_00025_));
 sky130_fd_sc_hd__o32a_1 _13499_ (.A1(_05485_),
    .A2(_08447_),
    .A3(_08520_),
    .B1(_08522_),
    .B2(net1581),
    .X(_00026_));
 sky130_fd_sc_hd__nand2_1 _13500_ (.A(_05886_),
    .B(_08443_),
    .Y(_08526_));
 sky130_fd_sc_hd__o32a_1 _13501_ (.A1(_05485_),
    .A2(_08526_),
    .A3(_08520_),
    .B1(_08522_),
    .B2(\min_sad_reg[12] ),
    .X(_00027_));
 sky130_fd_sc_hd__nand2_1 _13502_ (.A(_05886_),
    .B(_08440_),
    .Y(_08527_));
 sky130_fd_sc_hd__o32a_1 _13503_ (.A1(_05485_),
    .A2(_08527_),
    .A3(_08520_),
    .B1(_08522_),
    .B2(\min_sad_reg[13] ),
    .X(_00028_));
 sky130_fd_sc_hd__inv_2 _13504_ (.A(_08438_),
    .Y(_08528_));
 sky130_fd_sc_hd__o32a_1 _13505_ (.A1(_05485_),
    .A2(_08528_),
    .A3(_08520_),
    .B1(_08522_),
    .B2(\min_sad_reg[14] ),
    .X(_00029_));
 sky130_fd_sc_hd__nand2_1 _13506_ (.A(_05886_),
    .B(_08434_),
    .Y(_08529_));
 sky130_fd_sc_hd__o32a_1 _13507_ (.A1(_05485_),
    .A2(_08529_),
    .A3(_08520_),
    .B1(_08522_),
    .B2(net1962),
    .X(_00030_));
 sky130_fd_sc_hd__buf_12 _13508_ (.A(net97),
    .X(_08530_));
 sky130_fd_sc_hd__buf_8 _13509_ (.A(_08530_),
    .X(_08531_));
 sky130_fd_sc_hd__nand2_8 _13510_ (.A(net279),
    .B(\state[4] ),
    .Y(_08532_));
 sky130_fd_sc_hd__nor2_8 _13511_ (.A(_04433_),
    .B(_08532_),
    .Y(_08533_));
 sky130_fd_sc_hd__mux2_1 _13512_ (.A0(net1672),
    .A1(_08531_),
    .S(_08533_),
    .X(_08534_));
 sky130_fd_sc_hd__clkbuf_1 _13513_ (.A(_08534_),
    .X(_00031_));
 sky130_fd_sc_hd__clkbuf_8 _13514_ (.A(net98),
    .X(_08535_));
 sky130_fd_sc_hd__buf_6 _13515_ (.A(_08535_),
    .X(_08536_));
 sky130_fd_sc_hd__mux2_1 _13516_ (.A0(net699),
    .A1(_08536_),
    .S(_08533_),
    .X(_08537_));
 sky130_fd_sc_hd__clkbuf_1 _13517_ (.A(_08537_),
    .X(_00032_));
 sky130_fd_sc_hd__buf_8 _13518_ (.A(net99),
    .X(_08538_));
 sky130_fd_sc_hd__buf_8 _13519_ (.A(_08538_),
    .X(_08539_));
 sky130_fd_sc_hd__mux2_1 _13520_ (.A0(net1682),
    .A1(_08539_),
    .S(_08533_),
    .X(_08540_));
 sky130_fd_sc_hd__clkbuf_1 _13521_ (.A(_08540_),
    .X(_00033_));
 sky130_fd_sc_hd__buf_8 _13522_ (.A(net100),
    .X(_08541_));
 sky130_fd_sc_hd__clkbuf_16 _13523_ (.A(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__mux2_1 _13524_ (.A0(net1940),
    .A1(_08542_),
    .S(_08533_),
    .X(_08543_));
 sky130_fd_sc_hd__clkbuf_1 _13525_ (.A(_08543_),
    .X(_00034_));
 sky130_fd_sc_hd__buf_8 _13526_ (.A(net101),
    .X(_08544_));
 sky130_fd_sc_hd__clkbuf_16 _13527_ (.A(_08544_),
    .X(_08545_));
 sky130_fd_sc_hd__mux2_1 _13528_ (.A0(net725),
    .A1(_08545_),
    .S(_08533_),
    .X(_08546_));
 sky130_fd_sc_hd__clkbuf_1 _13529_ (.A(_08546_),
    .X(_00035_));
 sky130_fd_sc_hd__buf_8 _13530_ (.A(net102),
    .X(_08547_));
 sky130_fd_sc_hd__clkbuf_16 _13531_ (.A(_08547_),
    .X(_08548_));
 sky130_fd_sc_hd__mux2_1 _13532_ (.A0(net1113),
    .A1(_08548_),
    .S(_08533_),
    .X(_08549_));
 sky130_fd_sc_hd__clkbuf_1 _13533_ (.A(_08549_),
    .X(_00036_));
 sky130_fd_sc_hd__buf_4 _13534_ (.A(net103),
    .X(_08550_));
 sky130_fd_sc_hd__buf_6 _13535_ (.A(_08550_),
    .X(_08551_));
 sky130_fd_sc_hd__mux2_1 _13536_ (.A0(net677),
    .A1(_08551_),
    .S(_08533_),
    .X(_08552_));
 sky130_fd_sc_hd__clkbuf_1 _13537_ (.A(_08552_),
    .X(_00037_));
 sky130_fd_sc_hd__buf_4 _13538_ (.A(net104),
    .X(_08553_));
 sky130_fd_sc_hd__clkbuf_8 _13539_ (.A(_08553_),
    .X(_08554_));
 sky130_fd_sc_hd__mux2_1 _13540_ (.A0(net1250),
    .A1(_08554_),
    .S(_08533_),
    .X(_08555_));
 sky130_fd_sc_hd__clkbuf_1 _13541_ (.A(_08555_),
    .X(_00038_));
 sky130_fd_sc_hd__and2_1 _13542_ (.A(_04447_),
    .B(_04436_),
    .X(_08556_));
 sky130_fd_sc_hd__buf_4 _13543_ (.A(\state[6] ),
    .X(_08557_));
 sky130_fd_sc_hd__or2_1 _13544_ (.A(_04442_),
    .B(_08508_),
    .X(_08558_));
 sky130_fd_sc_hd__nand2_1 _13545_ (.A(_08557_),
    .B(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__o211a_1 _13546_ (.A1(_08557_),
    .A2(\state[2] ),
    .B1(_08559_),
    .C1(net272),
    .X(_08560_));
 sky130_fd_sc_hd__mux2_1 _13547_ (.A0(net727),
    .A1(_08556_),
    .S(_08560_),
    .X(_08561_));
 sky130_fd_sc_hd__clkbuf_1 _13548_ (.A(_08561_),
    .X(_00039_));
 sky130_fd_sc_hd__and2_1 _13549_ (.A(_04447_),
    .B(_04437_),
    .X(_08562_));
 sky130_fd_sc_hd__mux2_1 _13550_ (.A0(net599),
    .A1(_08562_),
    .S(_08560_),
    .X(_08563_));
 sky130_fd_sc_hd__clkbuf_1 _13551_ (.A(_08563_),
    .X(_00040_));
 sky130_fd_sc_hd__and2_1 _13552_ (.A(_04447_),
    .B(_04435_),
    .X(_08564_));
 sky130_fd_sc_hd__mux2_1 _13553_ (.A0(net291),
    .A1(_08564_),
    .S(_08560_),
    .X(_08565_));
 sky130_fd_sc_hd__clkbuf_1 _13554_ (.A(_08565_),
    .X(_00041_));
 sky130_fd_sc_hd__and2_1 _13555_ (.A(\point_cnt[3] ),
    .B(_04447_),
    .X(_08566_));
 sky130_fd_sc_hd__mux2_1 _13556_ (.A0(net398),
    .A1(_08566_),
    .S(_08560_),
    .X(_08567_));
 sky130_fd_sc_hd__clkbuf_1 _13557_ (.A(_08567_),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_1 _13558_ (.A0(net172),
    .A1(\best_cand_x[0] ),
    .S(_04449_),
    .X(_08568_));
 sky130_fd_sc_hd__clkbuf_1 _13559_ (.A(_08568_),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_1 _13560_ (.A0(net173),
    .A1(net1597),
    .S(_04449_),
    .X(_08569_));
 sky130_fd_sc_hd__clkbuf_1 _13561_ (.A(_08569_),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _13562_ (.A0(net174),
    .A1(net1839),
    .S(_04449_),
    .X(_08570_));
 sky130_fd_sc_hd__clkbuf_1 _13563_ (.A(_08570_),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _13564_ (.A0(net175),
    .A1(net1602),
    .S(_04449_),
    .X(_08571_));
 sky130_fd_sc_hd__clkbuf_1 _13565_ (.A(_08571_),
    .X(_00046_));
 sky130_fd_sc_hd__mux2_1 _13566_ (.A0(net176),
    .A1(net1787),
    .S(_04449_),
    .X(_08572_));
 sky130_fd_sc_hd__clkbuf_1 _13567_ (.A(_08572_),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _13568_ (.A0(net177),
    .A1(\best_cand_x[5] ),
    .S(_04449_),
    .X(_08573_));
 sky130_fd_sc_hd__clkbuf_1 _13569_ (.A(_08573_),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _13570_ (.A0(net178),
    .A1(net975),
    .S(_04449_),
    .X(_08574_));
 sky130_fd_sc_hd__clkbuf_1 _13571_ (.A(_08574_),
    .X(_00049_));
 sky130_fd_sc_hd__buf_6 _13572_ (.A(\state[7] ),
    .X(_08575_));
 sky130_fd_sc_hd__mux2_1 _13573_ (.A0(net179),
    .A1(net1998),
    .S(_08575_),
    .X(_08576_));
 sky130_fd_sc_hd__clkbuf_1 _13574_ (.A(_08576_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _13575_ (.A0(net180),
    .A1(\best_cand_y[2] ),
    .S(_08575_),
    .X(_08577_));
 sky130_fd_sc_hd__clkbuf_1 _13576_ (.A(_08577_),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _13577_ (.A0(net181),
    .A1(\best_cand_y[3] ),
    .S(_08575_),
    .X(_08578_));
 sky130_fd_sc_hd__clkbuf_1 _13578_ (.A(_08578_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _13579_ (.A0(net182),
    .A1(net1880),
    .S(_08575_),
    .X(_08579_));
 sky130_fd_sc_hd__clkbuf_1 _13580_ (.A(_08579_),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _13581_ (.A0(net183),
    .A1(\best_cand_y[5] ),
    .S(_08575_),
    .X(_08580_));
 sky130_fd_sc_hd__clkbuf_1 _13582_ (.A(_08580_),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _13583_ (.A0(net1938),
    .A1(\min_sad_reg[0] ),
    .S(_08575_),
    .X(_08581_));
 sky130_fd_sc_hd__clkbuf_1 _13584_ (.A(_08581_),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _13585_ (.A0(net191),
    .A1(\min_sad_reg[1] ),
    .S(_08575_),
    .X(_08582_));
 sky130_fd_sc_hd__clkbuf_1 _13586_ (.A(_08582_),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _13587_ (.A0(net192),
    .A1(\min_sad_reg[2] ),
    .S(_08575_),
    .X(_08583_));
 sky130_fd_sc_hd__clkbuf_1 _13588_ (.A(_08583_),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _13589_ (.A0(net1891),
    .A1(\min_sad_reg[3] ),
    .S(_08575_),
    .X(_08584_));
 sky130_fd_sc_hd__clkbuf_1 _13590_ (.A(_08584_),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _13591_ (.A0(net1819),
    .A1(\min_sad_reg[4] ),
    .S(_08575_),
    .X(_08585_));
 sky130_fd_sc_hd__clkbuf_1 _13592_ (.A(_08585_),
    .X(_00059_));
 sky130_fd_sc_hd__buf_8 _13593_ (.A(\state[7] ),
    .X(_08586_));
 sky130_fd_sc_hd__mux2_1 _13594_ (.A0(net195),
    .A1(\min_sad_reg[5] ),
    .S(_08586_),
    .X(_08587_));
 sky130_fd_sc_hd__clkbuf_1 _13595_ (.A(_08587_),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _13596_ (.A0(net196),
    .A1(\min_sad_reg[6] ),
    .S(_08586_),
    .X(_08588_));
 sky130_fd_sc_hd__clkbuf_1 _13597_ (.A(_08588_),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _13598_ (.A0(net1829),
    .A1(\min_sad_reg[7] ),
    .S(_08586_),
    .X(_08589_));
 sky130_fd_sc_hd__clkbuf_1 _13599_ (.A(_08589_),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _13600_ (.A0(net198),
    .A1(\min_sad_reg[8] ),
    .S(_08586_),
    .X(_08590_));
 sky130_fd_sc_hd__clkbuf_1 _13601_ (.A(_08590_),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _13602_ (.A0(net199),
    .A1(\min_sad_reg[9] ),
    .S(_08586_),
    .X(_08591_));
 sky130_fd_sc_hd__clkbuf_1 _13603_ (.A(_08591_),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _13604_ (.A0(net185),
    .A1(\min_sad_reg[10] ),
    .S(_08586_),
    .X(_08592_));
 sky130_fd_sc_hd__clkbuf_1 _13605_ (.A(_08592_),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _13606_ (.A0(net186),
    .A1(\min_sad_reg[11] ),
    .S(_08586_),
    .X(_08593_));
 sky130_fd_sc_hd__clkbuf_1 _13607_ (.A(_08593_),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _13608_ (.A0(net187),
    .A1(\min_sad_reg[12] ),
    .S(_08586_),
    .X(_08594_));
 sky130_fd_sc_hd__clkbuf_1 _13609_ (.A(_08594_),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _13610_ (.A0(net188),
    .A1(\min_sad_reg[13] ),
    .S(_08586_),
    .X(_08595_));
 sky130_fd_sc_hd__clkbuf_1 _13611_ (.A(_08595_),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _13612_ (.A0(net189),
    .A1(\min_sad_reg[14] ),
    .S(_08586_),
    .X(_08596_));
 sky130_fd_sc_hd__clkbuf_1 _13613_ (.A(_08596_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _13614_ (.A0(net190),
    .A1(\min_sad_reg[15] ),
    .S(\state[7] ),
    .X(_08597_));
 sky130_fd_sc_hd__clkbuf_1 _13615_ (.A(_08597_),
    .X(_00070_));
 sky130_fd_sc_hd__inv_2 _13616_ (.A(net1997),
    .Y(_08598_));
 sky130_fd_sc_hd__a21o_1 _13617_ (.A1(_08598_),
    .A2(net139),
    .B1(_04449_),
    .X(_00071_));
 sky130_fd_sc_hd__and2_1 _13618_ (.A(_04455_),
    .B(\best_cand_x[0] ),
    .X(_08599_));
 sky130_fd_sc_hd__nor2_1 _13619_ (.A(_04443_),
    .B(\state[1] ),
    .Y(_08600_));
 sky130_fd_sc_hd__a211o_2 _13620_ (.A1(_04443_),
    .A2(_04442_),
    .B1(_00002_),
    .C1(_08600_),
    .X(_08601_));
 sky130_fd_sc_hd__buf_4 _13621_ (.A(_08601_),
    .X(_08602_));
 sky130_fd_sc_hd__mux2_1 _13622_ (.A0(_08599_),
    .A1(\center_x[0] ),
    .S(_08602_),
    .X(_08603_));
 sky130_fd_sc_hd__clkbuf_1 _13623_ (.A(_08603_),
    .X(_00072_));
 sky130_fd_sc_hd__and2_1 _13624_ (.A(_04455_),
    .B(\best_cand_x[1] ),
    .X(_08604_));
 sky130_fd_sc_hd__mux2_1 _13625_ (.A0(_08604_),
    .A1(\center_x[1] ),
    .S(_08602_),
    .X(_08605_));
 sky130_fd_sc_hd__clkbuf_1 _13626_ (.A(_08605_),
    .X(_00073_));
 sky130_fd_sc_hd__and2_1 _13627_ (.A(_04455_),
    .B(\best_cand_x[2] ),
    .X(_08606_));
 sky130_fd_sc_hd__mux2_1 _13628_ (.A0(_08606_),
    .A1(\center_x[2] ),
    .S(_08602_),
    .X(_08607_));
 sky130_fd_sc_hd__clkbuf_1 _13629_ (.A(_08607_),
    .X(_00074_));
 sky130_fd_sc_hd__and2_1 _13630_ (.A(_04455_),
    .B(\best_cand_x[3] ),
    .X(_08608_));
 sky130_fd_sc_hd__mux2_1 _13631_ (.A0(_08608_),
    .A1(\center_x[3] ),
    .S(_08602_),
    .X(_08609_));
 sky130_fd_sc_hd__clkbuf_1 _13632_ (.A(_08609_),
    .X(_00075_));
 sky130_fd_sc_hd__and2_1 _13633_ (.A(_04455_),
    .B(\best_cand_x[4] ),
    .X(_08610_));
 sky130_fd_sc_hd__mux2_1 _13634_ (.A0(_08610_),
    .A1(\center_x[4] ),
    .S(_08602_),
    .X(_08611_));
 sky130_fd_sc_hd__clkbuf_1 _13635_ (.A(_08611_),
    .X(_00076_));
 sky130_fd_sc_hd__and2_1 _13636_ (.A(_04455_),
    .B(\best_cand_x[5] ),
    .X(_08612_));
 sky130_fd_sc_hd__mux2_1 _13637_ (.A0(_08612_),
    .A1(\center_x[5] ),
    .S(_08602_),
    .X(_08613_));
 sky130_fd_sc_hd__clkbuf_1 _13638_ (.A(_08613_),
    .X(_00077_));
 sky130_fd_sc_hd__and2_1 _13639_ (.A(_04455_),
    .B(\best_cand_x[6] ),
    .X(_08614_));
 sky130_fd_sc_hd__mux2_1 _13640_ (.A0(_08614_),
    .A1(\center_x[6] ),
    .S(_08602_),
    .X(_08615_));
 sky130_fd_sc_hd__clkbuf_1 _13641_ (.A(_08615_),
    .X(_00078_));
 sky130_fd_sc_hd__and2_1 _13642_ (.A(_04455_),
    .B(\best_cand_y[0] ),
    .X(_08616_));
 sky130_fd_sc_hd__mux2_1 _13643_ (.A0(_08616_),
    .A1(\center_y[0] ),
    .S(_08602_),
    .X(_08617_));
 sky130_fd_sc_hd__clkbuf_1 _13644_ (.A(_08617_),
    .X(_00079_));
 sky130_fd_sc_hd__inv_2 _13645_ (.A(\center_y[1] ),
    .Y(_08618_));
 sky130_fd_sc_hd__a21oi_1 _13646_ (.A1(_04455_),
    .A2(net1569),
    .B1(_08602_),
    .Y(_08619_));
 sky130_fd_sc_hd__a21oi_1 _13647_ (.A1(_08618_),
    .A2(_08602_),
    .B1(_08619_),
    .Y(_00080_));
 sky130_fd_sc_hd__and2_1 _13648_ (.A(\state[1] ),
    .B(\best_cand_y[2] ),
    .X(_08620_));
 sky130_fd_sc_hd__mux2_1 _13649_ (.A0(_08620_),
    .A1(\center_y[2] ),
    .S(_08601_),
    .X(_08621_));
 sky130_fd_sc_hd__clkbuf_1 _13650_ (.A(_08621_),
    .X(_00081_));
 sky130_fd_sc_hd__and2_1 _13651_ (.A(\state[1] ),
    .B(\best_cand_y[3] ),
    .X(_08622_));
 sky130_fd_sc_hd__mux2_1 _13652_ (.A0(_08622_),
    .A1(\center_y[3] ),
    .S(_08601_),
    .X(_08623_));
 sky130_fd_sc_hd__clkbuf_1 _13653_ (.A(_08623_),
    .X(_00082_));
 sky130_fd_sc_hd__and2_1 _13654_ (.A(\state[1] ),
    .B(\best_cand_y[4] ),
    .X(_08624_));
 sky130_fd_sc_hd__mux2_1 _13655_ (.A0(_08624_),
    .A1(\center_y[4] ),
    .S(_08601_),
    .X(_08625_));
 sky130_fd_sc_hd__clkbuf_1 _13656_ (.A(_08625_),
    .X(_00083_));
 sky130_fd_sc_hd__and2_1 _13657_ (.A(\state[1] ),
    .B(\best_cand_y[5] ),
    .X(_08626_));
 sky130_fd_sc_hd__mux2_1 _13658_ (.A0(_08626_),
    .A1(\center_y[5] ),
    .S(_08601_),
    .X(_08627_));
 sky130_fd_sc_hd__clkbuf_1 _13659_ (.A(_08627_),
    .X(_00084_));
 sky130_fd_sc_hd__and2_1 _13660_ (.A(\state[1] ),
    .B(\best_cand_y[6] ),
    .X(_08628_));
 sky130_fd_sc_hd__mux2_1 _13661_ (.A0(_08628_),
    .A1(\center_y[6] ),
    .S(_08601_),
    .X(_08629_));
 sky130_fd_sc_hd__clkbuf_1 _13662_ (.A(_08629_),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _13663_ (.A0(\center_x[0] ),
    .A1(\cand_x[0] ),
    .S(_04454_),
    .X(_08630_));
 sky130_fd_sc_hd__or2_2 _13664_ (.A(_04453_),
    .B(shex_load),
    .X(_08631_));
 sky130_fd_sc_hd__a2bb2o_2 _13665_ (.A1_N(_08558_),
    .A2_N(_08631_),
    .B1(\state[5] ),
    .B2(_04453_),
    .X(_08632_));
 sky130_fd_sc_hd__buf_4 _13666_ (.A(_08632_),
    .X(_08633_));
 sky130_fd_sc_hd__mux2_1 _13667_ (.A0(net1961),
    .A1(_08630_),
    .S(_08633_),
    .X(_08634_));
 sky130_fd_sc_hd__clkbuf_1 _13668_ (.A(_08634_),
    .X(_00086_));
 sky130_fd_sc_hd__buf_4 _13669_ (.A(\state[3] ),
    .X(_08635_));
 sky130_fd_sc_hd__mux2_1 _13670_ (.A0(\center_x[1] ),
    .A1(\cand_x[1] ),
    .S(_08635_),
    .X(_08636_));
 sky130_fd_sc_hd__mux2_1 _13671_ (.A0(\shex_center_x[1] ),
    .A1(_08636_),
    .S(_08633_),
    .X(_08637_));
 sky130_fd_sc_hd__clkbuf_1 _13672_ (.A(_08637_),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _13673_ (.A0(\center_x[2] ),
    .A1(\cand_x[2] ),
    .S(_08635_),
    .X(_08638_));
 sky130_fd_sc_hd__mux2_1 _13674_ (.A0(\shex_center_x[2] ),
    .A1(_08638_),
    .S(_08633_),
    .X(_08639_));
 sky130_fd_sc_hd__clkbuf_1 _13675_ (.A(_08639_),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _13676_ (.A0(\center_x[3] ),
    .A1(\cand_x[3] ),
    .S(_08635_),
    .X(_08640_));
 sky130_fd_sc_hd__mux2_1 _13677_ (.A0(net1921),
    .A1(_08640_),
    .S(_08633_),
    .X(_08641_));
 sky130_fd_sc_hd__clkbuf_1 _13678_ (.A(_08641_),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _13679_ (.A0(\center_x[4] ),
    .A1(\cand_x[4] ),
    .S(_08635_),
    .X(_08642_));
 sky130_fd_sc_hd__mux2_1 _13680_ (.A0(net1960),
    .A1(_08642_),
    .S(_08633_),
    .X(_08643_));
 sky130_fd_sc_hd__clkbuf_1 _13681_ (.A(_08643_),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _13682_ (.A0(\center_x[5] ),
    .A1(\cand_x[5] ),
    .S(_08635_),
    .X(_08644_));
 sky130_fd_sc_hd__mux2_1 _13683_ (.A0(net1952),
    .A1(_08644_),
    .S(_08633_),
    .X(_08645_));
 sky130_fd_sc_hd__clkbuf_1 _13684_ (.A(_08645_),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _13685_ (.A0(\center_x[6] ),
    .A1(_04475_),
    .S(_08635_),
    .X(_08646_));
 sky130_fd_sc_hd__mux2_1 _13686_ (.A0(net1929),
    .A1(_08646_),
    .S(_08633_),
    .X(_08647_));
 sky130_fd_sc_hd__clkbuf_1 _13687_ (.A(_08647_),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _13688_ (.A0(\center_y[0] ),
    .A1(\cand_y[0] ),
    .S(_08635_),
    .X(_08648_));
 sky130_fd_sc_hd__mux2_1 _13689_ (.A0(\shex_center_y[0] ),
    .A1(_08648_),
    .S(_08633_),
    .X(_08649_));
 sky130_fd_sc_hd__clkbuf_1 _13690_ (.A(_08649_),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _13691_ (.A0(\center_y[1] ),
    .A1(\cand_y[1] ),
    .S(_08635_),
    .X(_08650_));
 sky130_fd_sc_hd__mux2_1 _13692_ (.A0(net1916),
    .A1(_08650_),
    .S(_08633_),
    .X(_08651_));
 sky130_fd_sc_hd__clkbuf_1 _13693_ (.A(_08651_),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _13694_ (.A0(\center_y[2] ),
    .A1(\cand_y[2] ),
    .S(_08635_),
    .X(_08652_));
 sky130_fd_sc_hd__mux2_1 _13695_ (.A0(net1937),
    .A1(_08652_),
    .S(_08633_),
    .X(_08653_));
 sky130_fd_sc_hd__clkbuf_1 _13696_ (.A(_08653_),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _13697_ (.A0(\center_y[3] ),
    .A1(\cand_y[3] ),
    .S(_08635_),
    .X(_08654_));
 sky130_fd_sc_hd__mux2_1 _13698_ (.A0(net1948),
    .A1(_08654_),
    .S(_08632_),
    .X(_08655_));
 sky130_fd_sc_hd__clkbuf_1 _13699_ (.A(_08655_),
    .X(_00096_));
 sky130_fd_sc_hd__buf_4 _13700_ (.A(\state[3] ),
    .X(_08656_));
 sky130_fd_sc_hd__mux2_1 _13701_ (.A0(\center_y[4] ),
    .A1(\cand_y[4] ),
    .S(_08656_),
    .X(_08657_));
 sky130_fd_sc_hd__mux2_1 _13702_ (.A0(\shex_center_y[4] ),
    .A1(_08657_),
    .S(_08632_),
    .X(_08658_));
 sky130_fd_sc_hd__clkbuf_1 _13703_ (.A(_08658_),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _13704_ (.A0(\center_y[5] ),
    .A1(\cand_y[5] ),
    .S(_08656_),
    .X(_08659_));
 sky130_fd_sc_hd__mux2_1 _13705_ (.A0(\shex_center_y[5] ),
    .A1(_08659_),
    .S(_08632_),
    .X(_08660_));
 sky130_fd_sc_hd__clkbuf_1 _13706_ (.A(_08660_),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _13707_ (.A0(\center_y[6] ),
    .A1(_04851_),
    .S(_08656_),
    .X(_08661_));
 sky130_fd_sc_hd__mux2_1 _13708_ (.A0(net1971),
    .A1(_08661_),
    .S(_08632_),
    .X(_08662_));
 sky130_fd_sc_hd__clkbuf_1 _13709_ (.A(_08662_),
    .X(_00099_));
 sky130_fd_sc_hd__nand2_1 _13710_ (.A(_04436_),
    .B(\shex_center_x[0] ),
    .Y(_08663_));
 sky130_fd_sc_hd__or2_1 _13711_ (.A(_04436_),
    .B(\shex_center_x[0] ),
    .X(_08664_));
 sky130_fd_sc_hd__o21a_1 _13712_ (.A1(_08557_),
    .A2(_04453_),
    .B1(\center_x[0] ),
    .X(_08665_));
 sky130_fd_sc_hd__a31o_1 _13713_ (.A1(_04454_),
    .A2(_08663_),
    .A3(_08664_),
    .B1(_08665_),
    .X(_08666_));
 sky130_fd_sc_hd__or2_1 _13714_ (.A(_04442_),
    .B(_04440_),
    .X(_08667_));
 sky130_fd_sc_hd__nand2_1 _13715_ (.A(\state[6] ),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__o211a_2 _13716_ (.A1(\state[2] ),
    .A2(_04462_),
    .B1(_08631_),
    .C1(_08668_),
    .X(_08669_));
 sky130_fd_sc_hd__buf_4 _13717_ (.A(_08669_),
    .X(_08670_));
 sky130_fd_sc_hd__mux2_1 _13718_ (.A0(\cand_x[0] ),
    .A1(_08666_),
    .S(_08670_),
    .X(_08671_));
 sky130_fd_sc_hd__clkbuf_1 _13719_ (.A(_08671_),
    .X(_00100_));
 sky130_fd_sc_hd__or3_1 _13720_ (.A(\point_cnt[2] ),
    .B(_04437_),
    .C(\point_cnt[0] ),
    .X(_08672_));
 sky130_fd_sc_hd__and2_1 _13721_ (.A(_04450_),
    .B(_08672_),
    .X(_08673_));
 sky130_fd_sc_hd__or2_1 _13722_ (.A(\center_x[1] ),
    .B(_08673_),
    .X(_08674_));
 sky130_fd_sc_hd__nand2_1 _13723_ (.A(\center_x[1] ),
    .B(_08673_),
    .Y(_08675_));
 sky130_fd_sc_hd__and3_1 _13724_ (.A(\point_cnt[1] ),
    .B(\point_cnt[0] ),
    .C(\shex_center_x[1] ),
    .X(_08676_));
 sky130_fd_sc_hd__and2_1 _13725_ (.A(\point_cnt[1] ),
    .B(\point_cnt[0] ),
    .X(_08677_));
 sky130_fd_sc_hd__clkbuf_4 _13726_ (.A(_08677_),
    .X(_08678_));
 sky130_fd_sc_hd__nor2_1 _13727_ (.A(\shex_center_x[1] ),
    .B(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__o21ai_1 _13728_ (.A1(_08676_),
    .A2(_08679_),
    .B1(_08663_),
    .Y(_08680_));
 sky130_fd_sc_hd__or3_1 _13729_ (.A(_08663_),
    .B(_08676_),
    .C(_08679_),
    .X(_08681_));
 sky130_fd_sc_hd__a32o_1 _13730_ (.A1(_08656_),
    .A2(_08680_),
    .A3(_08681_),
    .B1(\center_x[1] ),
    .B2(_04686_),
    .X(_08682_));
 sky130_fd_sc_hd__a31o_1 _13731_ (.A1(_04447_),
    .A2(_08674_),
    .A3(_08675_),
    .B1(_08682_),
    .X(_08683_));
 sky130_fd_sc_hd__mux2_1 _13732_ (.A0(\cand_x[1] ),
    .A1(_08683_),
    .S(_08670_),
    .X(_08684_));
 sky130_fd_sc_hd__clkbuf_1 _13733_ (.A(_08684_),
    .X(_00101_));
 sky130_fd_sc_hd__xnor2_1 _13734_ (.A(\shex_center_x[2] ),
    .B(_08678_),
    .Y(_08685_));
 sky130_fd_sc_hd__and2b_1 _13735_ (.A_N(_08676_),
    .B(_08681_),
    .X(_08686_));
 sky130_fd_sc_hd__nand2_1 _13736_ (.A(_08685_),
    .B(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__or2_1 _13737_ (.A(_08685_),
    .B(_08686_),
    .X(_08688_));
 sky130_fd_sc_hd__and3_1 _13738_ (.A(_04435_),
    .B(\center_x[2] ),
    .C(_04450_),
    .X(_08689_));
 sky130_fd_sc_hd__and2_1 _13739_ (.A(_04435_),
    .B(_04450_),
    .X(_08690_));
 sky130_fd_sc_hd__buf_2 _13740_ (.A(_08690_),
    .X(_08691_));
 sky130_fd_sc_hd__nor2_1 _13741_ (.A(\center_x[2] ),
    .B(_08691_),
    .Y(_08692_));
 sky130_fd_sc_hd__o21ai_1 _13742_ (.A1(_08689_),
    .A2(_08692_),
    .B1(_08675_),
    .Y(_08693_));
 sky130_fd_sc_hd__or3_1 _13743_ (.A(_08675_),
    .B(_08689_),
    .C(_08692_),
    .X(_08694_));
 sky130_fd_sc_hd__a32o_1 _13744_ (.A1(_08557_),
    .A2(_08693_),
    .A3(_08694_),
    .B1(\center_x[2] ),
    .B2(_04686_),
    .X(_08695_));
 sky130_fd_sc_hd__a31o_1 _13745_ (.A1(_04454_),
    .A2(_08687_),
    .A3(_08688_),
    .B1(_08695_),
    .X(_08696_));
 sky130_fd_sc_hd__mux2_1 _13746_ (.A0(\cand_x[2] ),
    .A1(_08696_),
    .S(_08670_),
    .X(_08697_));
 sky130_fd_sc_hd__clkbuf_1 _13747_ (.A(_08697_),
    .X(_00102_));
 sky130_fd_sc_hd__and3_1 _13748_ (.A(_04437_),
    .B(_04436_),
    .C(\shex_center_x[3] ),
    .X(_08698_));
 sky130_fd_sc_hd__nor2_1 _13749_ (.A(\shex_center_x[3] ),
    .B(_08678_),
    .Y(_08699_));
 sky130_fd_sc_hd__a21bo_1 _13750_ (.A1(\shex_center_x[2] ),
    .A2(_08678_),
    .B1_N(_08688_),
    .X(_08700_));
 sky130_fd_sc_hd__or3b_1 _13751_ (.A(_08698_),
    .B(_08699_),
    .C_N(_08700_),
    .X(_08701_));
 sky130_fd_sc_hd__o21bai_1 _13752_ (.A1(_08698_),
    .A2(_08699_),
    .B1_N(_08700_),
    .Y(_08702_));
 sky130_fd_sc_hd__nand2_1 _13753_ (.A(\center_x[2] ),
    .B(_08691_),
    .Y(_08703_));
 sky130_fd_sc_hd__and3_1 _13754_ (.A(_04435_),
    .B(\center_x[3] ),
    .C(_04450_),
    .X(_08704_));
 sky130_fd_sc_hd__nor2_1 _13755_ (.A(\center_x[3] ),
    .B(_08691_),
    .Y(_08705_));
 sky130_fd_sc_hd__a211o_1 _13756_ (.A1(_08703_),
    .A2(_08694_),
    .B1(_08704_),
    .C1(_08705_),
    .X(_08706_));
 sky130_fd_sc_hd__o211ai_1 _13757_ (.A1(_08704_),
    .A2(_08705_),
    .B1(_08703_),
    .C1(_08694_),
    .Y(_08707_));
 sky130_fd_sc_hd__a32o_1 _13758_ (.A1(_08557_),
    .A2(_08706_),
    .A3(_08707_),
    .B1(\center_x[3] ),
    .B2(_04686_),
    .X(_08708_));
 sky130_fd_sc_hd__a31o_1 _13759_ (.A1(_04454_),
    .A2(_08701_),
    .A3(_08702_),
    .B1(_08708_),
    .X(_08709_));
 sky130_fd_sc_hd__mux2_1 _13760_ (.A0(\cand_x[3] ),
    .A1(_08709_),
    .S(_08670_),
    .X(_08710_));
 sky130_fd_sc_hd__clkbuf_1 _13761_ (.A(_08710_),
    .X(_00103_));
 sky130_fd_sc_hd__and2b_1 _13762_ (.A_N(_08699_),
    .B(_08700_),
    .X(_08711_));
 sky130_fd_sc_hd__nand2_1 _13763_ (.A(\shex_center_x[4] ),
    .B(_08678_),
    .Y(_08712_));
 sky130_fd_sc_hd__or2_1 _13764_ (.A(\shex_center_x[4] ),
    .B(_08678_),
    .X(_08713_));
 sky130_fd_sc_hd__o211a_1 _13765_ (.A1(_08698_),
    .A2(_08711_),
    .B1(_08712_),
    .C1(_08713_),
    .X(_08714_));
 sky130_fd_sc_hd__inv_2 _13766_ (.A(_08714_),
    .Y(_08715_));
 sky130_fd_sc_hd__a211o_1 _13767_ (.A1(_08712_),
    .A2(_08713_),
    .B1(_08698_),
    .C1(_08711_),
    .X(_08716_));
 sky130_fd_sc_hd__and3_1 _13768_ (.A(_04435_),
    .B(\center_x[4] ),
    .C(_04450_),
    .X(_08717_));
 sky130_fd_sc_hd__nor2_1 _13769_ (.A(\center_x[4] ),
    .B(_08691_),
    .Y(_08718_));
 sky130_fd_sc_hd__or2b_1 _13770_ (.A(_08704_),
    .B_N(_08706_),
    .X(_08719_));
 sky130_fd_sc_hd__or3b_1 _13771_ (.A(_08717_),
    .B(_08718_),
    .C_N(_08719_),
    .X(_08720_));
 sky130_fd_sc_hd__o21bai_1 _13772_ (.A1(_08717_),
    .A2(_08718_),
    .B1_N(_08719_),
    .Y(_08721_));
 sky130_fd_sc_hd__a32o_1 _13773_ (.A1(_08557_),
    .A2(_08720_),
    .A3(_08721_),
    .B1(\center_x[4] ),
    .B2(_04686_),
    .X(_08722_));
 sky130_fd_sc_hd__a31o_1 _13774_ (.A1(_04454_),
    .A2(_08715_),
    .A3(_08716_),
    .B1(_08722_),
    .X(_08723_));
 sky130_fd_sc_hd__mux2_1 _13775_ (.A0(\cand_x[4] ),
    .A1(_08723_),
    .S(_08670_),
    .X(_08724_));
 sky130_fd_sc_hd__clkbuf_1 _13776_ (.A(_08724_),
    .X(_00104_));
 sky130_fd_sc_hd__nand2_1 _13777_ (.A(\shex_center_x[5] ),
    .B(_08678_),
    .Y(_08725_));
 sky130_fd_sc_hd__or2_1 _13778_ (.A(\shex_center_x[5] ),
    .B(_08678_),
    .X(_08726_));
 sky130_fd_sc_hd__nand2_1 _13779_ (.A(_08725_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__and2_1 _13780_ (.A(_08712_),
    .B(_08715_),
    .X(_08728_));
 sky130_fd_sc_hd__o21ai_1 _13781_ (.A1(_08727_),
    .A2(_08728_),
    .B1(_04454_),
    .Y(_08729_));
 sky130_fd_sc_hd__a21oi_1 _13782_ (.A1(_08727_),
    .A2(_08728_),
    .B1(_08729_),
    .Y(_08730_));
 sky130_fd_sc_hd__and2b_1 _13783_ (.A_N(_08718_),
    .B(_08719_),
    .X(_08731_));
 sky130_fd_sc_hd__nand2_1 _13784_ (.A(\center_x[5] ),
    .B(_08691_),
    .Y(_08732_));
 sky130_fd_sc_hd__or2_1 _13785_ (.A(\center_x[5] ),
    .B(_08691_),
    .X(_08733_));
 sky130_fd_sc_hd__o211a_1 _13786_ (.A1(_08717_),
    .A2(_08731_),
    .B1(_08732_),
    .C1(_08733_),
    .X(_08734_));
 sky130_fd_sc_hd__a211o_1 _13787_ (.A1(_08732_),
    .A2(_08733_),
    .B1(_08717_),
    .C1(_08731_),
    .X(_08735_));
 sky130_fd_sc_hd__and3b_1 _13788_ (.A_N(_08734_),
    .B(_04447_),
    .C(_08735_),
    .X(_08736_));
 sky130_fd_sc_hd__a21bo_1 _13789_ (.A1(\center_x[5] ),
    .A2(_04688_),
    .B1_N(_08669_),
    .X(_08737_));
 sky130_fd_sc_hd__o32a_1 _13790_ (.A1(_08730_),
    .A2(_08736_),
    .A3(_08737_),
    .B1(_08670_),
    .B2(\cand_x[5] ),
    .X(_00105_));
 sky130_fd_sc_hd__a21o_1 _13791_ (.A1(\center_x[5] ),
    .A2(_08691_),
    .B1(_08734_),
    .X(_08738_));
 sky130_fd_sc_hd__xor2_1 _13792_ (.A(\center_x[6] ),
    .B(_08691_),
    .X(_08739_));
 sky130_fd_sc_hd__nand2_1 _13793_ (.A(_08738_),
    .B(_08739_),
    .Y(_08740_));
 sky130_fd_sc_hd__o21a_1 _13794_ (.A1(_08738_),
    .A2(_08739_),
    .B1(_08557_),
    .X(_08741_));
 sky130_fd_sc_hd__o211a_1 _13795_ (.A1(_08715_),
    .A2(_08727_),
    .B1(_08725_),
    .C1(_08712_),
    .X(_08742_));
 sky130_fd_sc_hd__xnor2_1 _13796_ (.A(\shex_center_x[6] ),
    .B(_08678_),
    .Y(_08743_));
 sky130_fd_sc_hd__o21ai_1 _13797_ (.A1(_08742_),
    .A2(_08743_),
    .B1(_08656_),
    .Y(_08744_));
 sky130_fd_sc_hd__a21oi_1 _13798_ (.A1(_08742_),
    .A2(_08743_),
    .B1(_08744_),
    .Y(_08745_));
 sky130_fd_sc_hd__a221o_1 _13799_ (.A1(\center_x[6] ),
    .A2(_04687_),
    .B1(_08740_),
    .B2(_08741_),
    .C1(_08745_),
    .X(_08746_));
 sky130_fd_sc_hd__mux2_1 _13800_ (.A0(_04475_),
    .A1(_08746_),
    .S(_08670_),
    .X(_08747_));
 sky130_fd_sc_hd__clkbuf_1 _13801_ (.A(_08747_),
    .X(_00106_));
 sky130_fd_sc_hd__or2b_1 _13802_ (.A(\shex_center_y[0] ),
    .B_N(_04436_),
    .X(_08748_));
 sky130_fd_sc_hd__or2b_1 _13803_ (.A(_04436_),
    .B_N(\shex_center_y[0] ),
    .X(_08749_));
 sky130_fd_sc_hd__and3_1 _13804_ (.A(\center_y[0] ),
    .B(_04450_),
    .C(_08672_),
    .X(_08750_));
 sky130_fd_sc_hd__o21ai_1 _13805_ (.A1(\center_y[0] ),
    .A2(_08673_),
    .B1(\state[6] ),
    .Y(_08751_));
 sky130_fd_sc_hd__a2bb2o_1 _13806_ (.A1_N(_08750_),
    .A2_N(_08751_),
    .B1(\center_y[0] ),
    .B2(_04686_),
    .X(_08752_));
 sky130_fd_sc_hd__a31o_1 _13807_ (.A1(_04454_),
    .A2(_08748_),
    .A3(_08749_),
    .B1(_08752_),
    .X(_08753_));
 sky130_fd_sc_hd__mux2_1 _13808_ (.A0(\cand_y[0] ),
    .A1(_08753_),
    .S(_08670_),
    .X(_08754_));
 sky130_fd_sc_hd__clkbuf_1 _13809_ (.A(_08754_),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _13810_ (.A0(_04436_),
    .A1(\point_cnt[2] ),
    .S(_04437_),
    .X(_08755_));
 sky130_fd_sc_hd__nor2_1 _13811_ (.A(_08618_),
    .B(_08755_),
    .Y(_08756_));
 sky130_fd_sc_hd__and2_1 _13812_ (.A(_08618_),
    .B(_08755_),
    .X(_08757_));
 sky130_fd_sc_hd__nor2_1 _13813_ (.A(_08756_),
    .B(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__xor2_1 _13814_ (.A(_08750_),
    .B(_08758_),
    .X(_08759_));
 sky130_fd_sc_hd__nor2_1 _13815_ (.A(\shex_center_y[1] ),
    .B(_04438_),
    .Y(_08760_));
 sky130_fd_sc_hd__and2_1 _13816_ (.A(\shex_center_y[1] ),
    .B(_04438_),
    .X(_08761_));
 sky130_fd_sc_hd__o21ai_1 _13817_ (.A1(_08760_),
    .A2(_08761_),
    .B1(_08749_),
    .Y(_08762_));
 sky130_fd_sc_hd__o311a_1 _13818_ (.A1(_08749_),
    .A2(_08760_),
    .A3(_08761_),
    .B1(_08762_),
    .C1(_08656_),
    .X(_08763_));
 sky130_fd_sc_hd__a221o_1 _13819_ (.A1(\center_y[1] ),
    .A2(_04687_),
    .B1(_08759_),
    .B2(_04447_),
    .C1(_08763_),
    .X(_08764_));
 sky130_fd_sc_hd__mux2_1 _13820_ (.A0(\cand_y[1] ),
    .A1(_08764_),
    .S(_08670_),
    .X(_08765_));
 sky130_fd_sc_hd__clkbuf_1 _13821_ (.A(_08765_),
    .X(_00108_));
 sky130_fd_sc_hd__o21ba_1 _13822_ (.A1(_04435_),
    .A2(_04437_),
    .B1_N(_08755_),
    .X(_08766_));
 sky130_fd_sc_hd__clkbuf_4 _13823_ (.A(_08766_),
    .X(_08767_));
 sky130_fd_sc_hd__xnor2_1 _13824_ (.A(\center_y[2] ),
    .B(_08767_),
    .Y(_08768_));
 sky130_fd_sc_hd__a21oi_1 _13825_ (.A1(_08750_),
    .A2(_08758_),
    .B1(_08756_),
    .Y(_08769_));
 sky130_fd_sc_hd__nand2_1 _13826_ (.A(_08768_),
    .B(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__or2_1 _13827_ (.A(_08768_),
    .B(_08769_),
    .X(_08771_));
 sky130_fd_sc_hd__or2_1 _13828_ (.A(\shex_center_y[2] ),
    .B(_04439_),
    .X(_08772_));
 sky130_fd_sc_hd__nand2_1 _13829_ (.A(\shex_center_y[2] ),
    .B(_04439_),
    .Y(_08773_));
 sky130_fd_sc_hd__nand2_1 _13830_ (.A(_08772_),
    .B(_08773_),
    .Y(_08774_));
 sky130_fd_sc_hd__o21ba_1 _13831_ (.A1(_08749_),
    .A2(_08760_),
    .B1_N(_08761_),
    .X(_08775_));
 sky130_fd_sc_hd__nand2_1 _13832_ (.A(_08774_),
    .B(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__or2_1 _13833_ (.A(_08774_),
    .B(_08775_),
    .X(_08777_));
 sky130_fd_sc_hd__a32o_1 _13834_ (.A1(_08656_),
    .A2(_08776_),
    .A3(_08777_),
    .B1(\center_y[2] ),
    .B2(_04686_),
    .X(_08778_));
 sky130_fd_sc_hd__a31o_1 _13835_ (.A1(_04447_),
    .A2(_08770_),
    .A3(_08771_),
    .B1(_08778_),
    .X(_08779_));
 sky130_fd_sc_hd__mux2_1 _13836_ (.A0(\cand_y[2] ),
    .A1(_08779_),
    .S(_08669_),
    .X(_08780_));
 sky130_fd_sc_hd__clkbuf_1 _13837_ (.A(_08780_),
    .X(_00109_));
 sky130_fd_sc_hd__a21bo_1 _13838_ (.A1(\center_y[2] ),
    .A2(_08767_),
    .B1_N(_08771_),
    .X(_08781_));
 sky130_fd_sc_hd__xnor2_1 _13839_ (.A(\center_y[3] ),
    .B(_08767_),
    .Y(_08782_));
 sky130_fd_sc_hd__xnor2_1 _13840_ (.A(_08781_),
    .B(_08782_),
    .Y(_08783_));
 sky130_fd_sc_hd__nor2_1 _13841_ (.A(\shex_center_y[3] ),
    .B(_04439_),
    .Y(_08784_));
 sky130_fd_sc_hd__nand2_1 _13842_ (.A(\shex_center_y[3] ),
    .B(_04439_),
    .Y(_08785_));
 sky130_fd_sc_hd__or2b_1 _13843_ (.A(_08784_),
    .B_N(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__and2_1 _13844_ (.A(_08773_),
    .B(_08777_),
    .X(_08787_));
 sky130_fd_sc_hd__o21ai_1 _13845_ (.A1(_08786_),
    .A2(_08787_),
    .B1(_08656_),
    .Y(_08788_));
 sky130_fd_sc_hd__a21oi_1 _13846_ (.A1(_08786_),
    .A2(_08787_),
    .B1(_08788_),
    .Y(_08789_));
 sky130_fd_sc_hd__a221o_1 _13847_ (.A1(\center_y[3] ),
    .A2(_04687_),
    .B1(_08783_),
    .B2(_08557_),
    .C1(_08789_),
    .X(_08790_));
 sky130_fd_sc_hd__mux2_1 _13848_ (.A0(\cand_y[3] ),
    .A1(_08790_),
    .S(_08669_),
    .X(_08791_));
 sky130_fd_sc_hd__clkbuf_1 _13849_ (.A(_08791_),
    .X(_00110_));
 sky130_fd_sc_hd__xnor2_1 _13850_ (.A(\center_y[4] ),
    .B(_08767_),
    .Y(_08792_));
 sky130_fd_sc_hd__o21ai_1 _13851_ (.A1(\center_y[2] ),
    .A2(\center_y[3] ),
    .B1(_08767_),
    .Y(_08793_));
 sky130_fd_sc_hd__o21a_1 _13852_ (.A1(_08771_),
    .A2(_08782_),
    .B1(_08793_),
    .X(_08794_));
 sky130_fd_sc_hd__nand2_1 _13853_ (.A(_08792_),
    .B(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__or2_1 _13854_ (.A(_08792_),
    .B(_08794_),
    .X(_08796_));
 sky130_fd_sc_hd__and3_1 _13855_ (.A(_04447_),
    .B(_08795_),
    .C(_08796_),
    .X(_08797_));
 sky130_fd_sc_hd__nor2_1 _13856_ (.A(\shex_center_y[4] ),
    .B(_04439_),
    .Y(_08798_));
 sky130_fd_sc_hd__and2_1 _13857_ (.A(\shex_center_y[4] ),
    .B(_04439_),
    .X(_08799_));
 sky130_fd_sc_hd__o21a_1 _13858_ (.A1(_08784_),
    .A2(_08787_),
    .B1(_08785_),
    .X(_08800_));
 sky130_fd_sc_hd__o21a_1 _13859_ (.A1(_08798_),
    .A2(_08799_),
    .B1(_08800_),
    .X(_08801_));
 sky130_fd_sc_hd__or3_1 _13860_ (.A(_08798_),
    .B(_08799_),
    .C(_08800_),
    .X(_08802_));
 sky130_fd_sc_hd__and3b_1 _13861_ (.A_N(_08801_),
    .B(_08802_),
    .C(_04454_),
    .X(_08803_));
 sky130_fd_sc_hd__a21bo_1 _13862_ (.A1(\center_y[4] ),
    .A2(_04688_),
    .B1_N(_08669_),
    .X(_08804_));
 sky130_fd_sc_hd__o32a_1 _13863_ (.A1(_08797_),
    .A2(_08803_),
    .A3(_08804_),
    .B1(_08670_),
    .B2(net306),
    .X(_00111_));
 sky130_fd_sc_hd__nand2_1 _13864_ (.A(\center_y[5] ),
    .B(_08767_),
    .Y(_08805_));
 sky130_fd_sc_hd__or2_1 _13865_ (.A(\center_y[5] ),
    .B(_08767_),
    .X(_08806_));
 sky130_fd_sc_hd__nand2_1 _13866_ (.A(_08805_),
    .B(_08806_),
    .Y(_08807_));
 sky130_fd_sc_hd__a21boi_1 _13867_ (.A1(\center_y[4] ),
    .A2(_08767_),
    .B1_N(_08796_),
    .Y(_08808_));
 sky130_fd_sc_hd__xor2_1 _13868_ (.A(_08807_),
    .B(_08808_),
    .X(_08809_));
 sky130_fd_sc_hd__xnor2_1 _13869_ (.A(\shex_center_y[5] ),
    .B(_04439_),
    .Y(_08810_));
 sky130_fd_sc_hd__and2b_1 _13870_ (.A_N(_08799_),
    .B(_08802_),
    .X(_08811_));
 sky130_fd_sc_hd__o21ai_1 _13871_ (.A1(_08810_),
    .A2(_08811_),
    .B1(_08656_),
    .Y(_08812_));
 sky130_fd_sc_hd__a21oi_1 _13872_ (.A1(_08810_),
    .A2(_08811_),
    .B1(_08812_),
    .Y(_08813_));
 sky130_fd_sc_hd__a221o_1 _13873_ (.A1(\center_y[5] ),
    .A2(_04687_),
    .B1(_08809_),
    .B2(_08557_),
    .C1(_08813_),
    .X(_08814_));
 sky130_fd_sc_hd__mux2_1 _13874_ (.A0(\cand_y[5] ),
    .A1(_08814_),
    .S(_08669_),
    .X(_08815_));
 sky130_fd_sc_hd__clkbuf_1 _13875_ (.A(_08815_),
    .X(_00112_));
 sky130_fd_sc_hd__nor2_1 _13876_ (.A(\center_y[5] ),
    .B(_08767_),
    .Y(_08816_));
 sky130_fd_sc_hd__o21ai_1 _13877_ (.A1(_08816_),
    .A2(_08808_),
    .B1(_08805_),
    .Y(_08817_));
 sky130_fd_sc_hd__xnor2_1 _13878_ (.A(\center_y[6] ),
    .B(_08767_),
    .Y(_08818_));
 sky130_fd_sc_hd__xnor2_1 _13879_ (.A(_08817_),
    .B(_08818_),
    .Y(_08819_));
 sky130_fd_sc_hd__o21ai_1 _13880_ (.A1(\shex_center_y[4] ),
    .A2(\shex_center_y[5] ),
    .B1(_04439_),
    .Y(_08820_));
 sky130_fd_sc_hd__o21a_1 _13881_ (.A1(_08802_),
    .A2(_08810_),
    .B1(_08820_),
    .X(_08821_));
 sky130_fd_sc_hd__xnor2_1 _13882_ (.A(\shex_center_y[6] ),
    .B(_04439_),
    .Y(_08822_));
 sky130_fd_sc_hd__o21ai_1 _13883_ (.A1(_08821_),
    .A2(_08822_),
    .B1(_08656_),
    .Y(_08823_));
 sky130_fd_sc_hd__a21oi_1 _13884_ (.A1(_08821_),
    .A2(_08822_),
    .B1(_08823_),
    .Y(_08824_));
 sky130_fd_sc_hd__a221o_1 _13885_ (.A1(\center_y[6] ),
    .A2(_04687_),
    .B1(_08819_),
    .B2(_08557_),
    .C1(_08824_),
    .X(_08825_));
 sky130_fd_sc_hd__mux2_1 _13886_ (.A0(_04851_),
    .A1(_08825_),
    .S(_08669_),
    .X(_08826_));
 sky130_fd_sc_hd__clkbuf_1 _13887_ (.A(_08826_),
    .X(_00113_));
 sky130_fd_sc_hd__nor2_1 _13888_ (.A(_04453_),
    .B(shex_load),
    .Y(_08827_));
 sky130_fd_sc_hd__or4_1 _13889_ (.A(\state[4] ),
    .B(\state[5] ),
    .C(\state[2] ),
    .D(_04462_),
    .X(_08828_));
 sky130_fd_sc_hd__mux2_1 _13890_ (.A0(net138),
    .A1(_08828_),
    .S(_08598_),
    .X(_08829_));
 sky130_fd_sc_hd__inv_2 _13891_ (.A(_08829_),
    .Y(_08830_));
 sky130_fd_sc_hd__a211o_4 _13892_ (.A1(_04434_),
    .A2(_08827_),
    .B1(_08830_),
    .C1(_00001_),
    .X(_08831_));
 sky130_fd_sc_hd__and3b_2 _13893_ (.A_N(\state[6] ),
    .B(_04955_),
    .C(_08631_),
    .X(_08832_));
 sky130_fd_sc_hd__nor2_2 _13894_ (.A(_08831_),
    .B(_08832_),
    .Y(_08833_));
 sky130_fd_sc_hd__mux2_1 _13895_ (.A0(_08833_),
    .A1(_08831_),
    .S(_04459_),
    .X(_08834_));
 sky130_fd_sc_hd__clkbuf_1 _13896_ (.A(_08834_),
    .X(_00114_));
 sky130_fd_sc_hd__nand2_1 _13897_ (.A(_04654_),
    .B(_04459_),
    .Y(_08835_));
 sky130_fd_sc_hd__a32o_1 _13898_ (.A1(_05887_),
    .A2(_08835_),
    .A3(_08833_),
    .B1(_08831_),
    .B2(_04654_),
    .X(_00115_));
 sky130_fd_sc_hd__nor2_1 _13899_ (.A(_08835_),
    .B(_08831_),
    .Y(_08836_));
 sky130_fd_sc_hd__a21oi_1 _13900_ (.A1(_04670_),
    .A2(_05898_),
    .B1(_08832_),
    .Y(_08837_));
 sky130_fd_sc_hd__or2_1 _13901_ (.A(_08831_),
    .B(_08837_),
    .X(_08838_));
 sky130_fd_sc_hd__o21a_1 _13902_ (.A1(_04670_),
    .A2(_08836_),
    .B1(_08838_),
    .X(_00116_));
 sky130_fd_sc_hd__buf_8 _13903_ (.A(_06103_),
    .X(_08839_));
 sky130_fd_sc_hd__a22o_1 _13904_ (.A1(_08839_),
    .A2(_08833_),
    .B1(_08838_),
    .B2(_04692_),
    .X(_00117_));
 sky130_fd_sc_hd__nor2_1 _13905_ (.A(_06176_),
    .B(_08831_),
    .Y(_08840_));
 sky130_fd_sc_hd__or3_4 _13906_ (.A(\state[6] ),
    .B(_04443_),
    .C(_08827_),
    .X(_08841_));
 sky130_fd_sc_hd__nand2_1 _13907_ (.A(_04738_),
    .B(_04424_),
    .Y(_08842_));
 sky130_fd_sc_hd__a21o_1 _13908_ (.A1(_08841_),
    .A2(_08842_),
    .B1(_08831_),
    .X(_08843_));
 sky130_fd_sc_hd__o21a_1 _13909_ (.A1(_04738_),
    .A2(_08840_),
    .B1(_08843_),
    .X(_00118_));
 sky130_fd_sc_hd__a32o_1 _13910_ (.A1(_04969_),
    .A2(_08841_),
    .A3(_08840_),
    .B1(_08843_),
    .B2(_04968_),
    .X(_00119_));
 sky130_fd_sc_hd__or2_1 _13911_ (.A(_05011_),
    .B(_08842_),
    .X(_08844_));
 sky130_fd_sc_hd__a21o_1 _13912_ (.A1(_08841_),
    .A2(_08844_),
    .B1(_08831_),
    .X(_08845_));
 sky130_fd_sc_hd__a21o_1 _13913_ (.A1(_05009_),
    .A2(_08840_),
    .B1(_05010_),
    .X(_08846_));
 sky130_fd_sc_hd__and2_1 _13914_ (.A(_08845_),
    .B(_08846_),
    .X(_08847_));
 sky130_fd_sc_hd__clkbuf_1 _13915_ (.A(_08847_),
    .X(_00120_));
 sky130_fd_sc_hd__a22o_1 _13916_ (.A1(_06101_),
    .A2(_08833_),
    .B1(_08845_),
    .B2(_05061_),
    .X(_00121_));
 sky130_fd_sc_hd__nor2_1 _13917_ (.A(_06304_),
    .B(_08832_),
    .Y(_08848_));
 sky130_fd_sc_hd__o21a_1 _13918_ (.A1(_08831_),
    .A2(_08848_),
    .B1(net297),
    .X(_00122_));
 sky130_fd_sc_hd__o31a_1 _13919_ (.A1(shex_load),
    .A2(_04442_),
    .A3(_04451_),
    .B1(\state[3] ),
    .X(_08849_));
 sky130_fd_sc_hd__a21oi_1 _13920_ (.A1(\state[6] ),
    .A2(_08667_),
    .B1(_08849_),
    .Y(_08850_));
 sky130_fd_sc_hd__or3_2 _13921_ (.A(\state[5] ),
    .B(\state[2] ),
    .C(_04462_),
    .X(_08851_));
 sky130_fd_sc_hd__a21o_1 _13922_ (.A1(_08850_),
    .A2(_08851_),
    .B1(_04436_),
    .X(_08852_));
 sky130_fd_sc_hd__o21ai_2 _13923_ (.A1(\state[5] ),
    .A2(\state[2] ),
    .B1(_08850_),
    .Y(_08853_));
 sky130_fd_sc_hd__and3_1 _13924_ (.A(_04436_),
    .B(_08850_),
    .C(_08851_),
    .X(_08854_));
 sky130_fd_sc_hd__inv_2 _13925_ (.A(_08854_),
    .Y(_08855_));
 sky130_fd_sc_hd__and3_1 _13926_ (.A(_08852_),
    .B(_08853_),
    .C(_08855_),
    .X(_08856_));
 sky130_fd_sc_hd__clkbuf_1 _13927_ (.A(_08856_),
    .X(_00123_));
 sky130_fd_sc_hd__or2_1 _13928_ (.A(_04437_),
    .B(_08854_),
    .X(_08857_));
 sky130_fd_sc_hd__and2_1 _13929_ (.A(_04437_),
    .B(_08854_),
    .X(_08858_));
 sky130_fd_sc_hd__inv_2 _13930_ (.A(_08858_),
    .Y(_08859_));
 sky130_fd_sc_hd__and3_1 _13931_ (.A(_08853_),
    .B(_08857_),
    .C(_08859_),
    .X(_08860_));
 sky130_fd_sc_hd__clkbuf_1 _13932_ (.A(_08860_),
    .X(_00124_));
 sky130_fd_sc_hd__or2_1 _13933_ (.A(_04435_),
    .B(_08858_),
    .X(_08861_));
 sky130_fd_sc_hd__and3_1 _13934_ (.A(_04435_),
    .B(_04437_),
    .C(_08854_),
    .X(_08862_));
 sky130_fd_sc_hd__inv_2 _13935_ (.A(_08862_),
    .Y(_08863_));
 sky130_fd_sc_hd__and3_1 _13936_ (.A(_08853_),
    .B(_08861_),
    .C(_08863_),
    .X(_08864_));
 sky130_fd_sc_hd__clkbuf_1 _13937_ (.A(_08864_),
    .X(_00125_));
 sky130_fd_sc_hd__o21ai_1 _13938_ (.A1(net309),
    .A2(_08862_),
    .B1(_08853_),
    .Y(_08865_));
 sky130_fd_sc_hd__a21oi_1 _13939_ (.A1(net309),
    .A2(_08862_),
    .B1(_08865_),
    .Y(_00126_));
 sky130_fd_sc_hd__nor3_1 _13940_ (.A(net310),
    .B(_04454_),
    .C(net1969),
    .Y(_08866_));
 sky130_fd_sc_hd__nor2_1 _13941_ (.A(_08849_),
    .B(_08866_),
    .Y(_00127_));
 sky130_fd_sc_hd__nand2_4 _13942_ (.A(net270),
    .B(_08851_),
    .Y(_08867_));
 sky130_fd_sc_hd__clkbuf_4 _13943_ (.A(_08867_),
    .X(_08868_));
 sky130_fd_sc_hd__or4b_2 _13944_ (.A(\state[5] ),
    .B(\state[3] ),
    .C(\state[2] ),
    .D_N(_08667_),
    .X(_08869_));
 sky130_fd_sc_hd__a21oi_4 _13945_ (.A1(_08631_),
    .A2(_08869_),
    .B1(_08867_),
    .Y(_08870_));
 sky130_fd_sc_hd__clkbuf_4 _13946_ (.A(_08870_),
    .X(_08871_));
 sky130_fd_sc_hd__a22o_1 _13947_ (.A1(net300),
    .A2(_08868_),
    .B1(_08871_),
    .B2(_08519_),
    .X(_00128_));
 sky130_fd_sc_hd__a22o_1 _13948_ (.A1(net301),
    .A2(_08868_),
    .B1(_08871_),
    .B2(_08478_),
    .X(_00129_));
 sky130_fd_sc_hd__a22o_1 _13949_ (.A1(net305),
    .A2(_08868_),
    .B1(_08871_),
    .B2(_08475_),
    .X(_00130_));
 sky130_fd_sc_hd__a22o_1 _13950_ (.A1(net295),
    .A2(_08868_),
    .B1(_08871_),
    .B2(_08488_),
    .X(_00131_));
 sky130_fd_sc_hd__a22o_1 _13951_ (.A1(net294),
    .A2(_08868_),
    .B1(_08871_),
    .B2(_08471_),
    .X(_00132_));
 sky130_fd_sc_hd__a22o_1 _13952_ (.A1(net293),
    .A2(_08868_),
    .B1(_08871_),
    .B2(_08524_),
    .X(_00133_));
 sky130_fd_sc_hd__a22o_1 _13953_ (.A1(net298),
    .A2(_08868_),
    .B1(_08871_),
    .B2(_08463_),
    .X(_00134_));
 sky130_fd_sc_hd__a22o_1 _13954_ (.A1(net304),
    .A2(_08868_),
    .B1(_08871_),
    .B2(_08461_),
    .X(_00135_));
 sky130_fd_sc_hd__a22o_1 _13955_ (.A1(net1638),
    .A2(_08868_),
    .B1(_08871_),
    .B2(_08456_),
    .X(_00136_));
 sky130_fd_sc_hd__a22o_1 _13956_ (.A1(net307),
    .A2(_08868_),
    .B1(_08871_),
    .B2(_08452_),
    .X(_00137_));
 sky130_fd_sc_hd__a22o_1 _13957_ (.A1(net308),
    .A2(_08867_),
    .B1(_08870_),
    .B2(_08525_),
    .X(_00138_));
 sky130_fd_sc_hd__a22o_1 _13958_ (.A1(net623),
    .A2(_08867_),
    .B1(_08870_),
    .B2(_08447_),
    .X(_00139_));
 sky130_fd_sc_hd__a22o_1 _13959_ (.A1(net303),
    .A2(_08867_),
    .B1(_08870_),
    .B2(_08526_),
    .X(_00140_));
 sky130_fd_sc_hd__a22o_1 _13960_ (.A1(net302),
    .A2(_08867_),
    .B1(_08870_),
    .B2(_08527_),
    .X(_00141_));
 sky130_fd_sc_hd__a22o_1 _13961_ (.A1(net299),
    .A2(_08867_),
    .B1(_08870_),
    .B2(_08528_),
    .X(_00142_));
 sky130_fd_sc_hd__a22o_1 _13962_ (.A1(net296),
    .A2(_08867_),
    .B1(_08870_),
    .B2(_08529_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _13963_ (.A0(\cand_y[0] ),
    .A1(net975),
    .S(_08511_),
    .X(_08872_));
 sky130_fd_sc_hd__clkbuf_1 _13964_ (.A(_08872_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _13965_ (.A0(\cand_y[1] ),
    .A1(net1999),
    .S(_08511_),
    .X(_08873_));
 sky130_fd_sc_hd__clkbuf_1 _13966_ (.A(_08873_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _13967_ (.A0(\cand_y[2] ),
    .A1(\best_cand_y[2] ),
    .S(_08511_),
    .X(_08874_));
 sky130_fd_sc_hd__clkbuf_1 _13968_ (.A(_08874_),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _13969_ (.A0(\cand_y[3] ),
    .A1(\best_cand_y[3] ),
    .S(_08510_),
    .X(_08875_));
 sky130_fd_sc_hd__clkbuf_1 _13970_ (.A(_08875_),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _13971_ (.A0(net306),
    .A1(net1880),
    .S(_08510_),
    .X(_08876_));
 sky130_fd_sc_hd__clkbuf_1 _13972_ (.A(_08876_),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _13973_ (.A0(\cand_y[5] ),
    .A1(\best_cand_y[5] ),
    .S(_08510_),
    .X(_08877_));
 sky130_fd_sc_hd__clkbuf_1 _13974_ (.A(_08877_),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _13975_ (.A0(_04851_),
    .A1(net698),
    .S(_08510_),
    .X(_08878_));
 sky130_fd_sc_hd__clkbuf_1 _13976_ (.A(_08878_),
    .X(_00150_));
 sky130_fd_sc_hd__clkbuf_16 _13977_ (.A(_08530_),
    .X(_08879_));
 sky130_fd_sc_hd__and2_4 _13978_ (.A(net280),
    .B(\state[4] ),
    .X(_08880_));
 sky130_fd_sc_hd__and2_1 _13979_ (.A(_05973_),
    .B(_08880_),
    .X(_08881_));
 sky130_fd_sc_hd__buf_12 _13980_ (.A(_08881_),
    .X(_08882_));
 sky130_fd_sc_hd__buf_12 _13981_ (.A(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__nand2_4 _13982_ (.A(_06113_),
    .B(_08883_),
    .Y(_08884_));
 sky130_fd_sc_hd__mux2_1 _13983_ (.A0(_08879_),
    .A1(\cur_mb_mem[0][0] ),
    .S(_08884_),
    .X(_08885_));
 sky130_fd_sc_hd__clkbuf_1 _13984_ (.A(_08885_),
    .X(_00151_));
 sky130_fd_sc_hd__buf_8 _13985_ (.A(_08535_),
    .X(_08886_));
 sky130_fd_sc_hd__mux2_1 _13986_ (.A0(_08886_),
    .A1(\cur_mb_mem[0][1] ),
    .S(_08884_),
    .X(_08887_));
 sky130_fd_sc_hd__clkbuf_1 _13987_ (.A(_08887_),
    .X(_00152_));
 sky130_fd_sc_hd__clkbuf_16 _13988_ (.A(_08538_),
    .X(_08888_));
 sky130_fd_sc_hd__mux2_1 _13989_ (.A0(_08888_),
    .A1(net1216),
    .S(_08884_),
    .X(_08889_));
 sky130_fd_sc_hd__clkbuf_1 _13990_ (.A(_08889_),
    .X(_00153_));
 sky130_fd_sc_hd__clkbuf_16 _13991_ (.A(_08541_),
    .X(_08890_));
 sky130_fd_sc_hd__mux2_1 _13992_ (.A0(_08890_),
    .A1(\cur_mb_mem[0][3] ),
    .S(_08884_),
    .X(_08891_));
 sky130_fd_sc_hd__clkbuf_1 _13993_ (.A(_08891_),
    .X(_00154_));
 sky130_fd_sc_hd__buf_8 _13994_ (.A(_08544_),
    .X(_08892_));
 sky130_fd_sc_hd__mux2_1 _13995_ (.A0(_08892_),
    .A1(\cur_mb_mem[0][4] ),
    .S(_08884_),
    .X(_08893_));
 sky130_fd_sc_hd__clkbuf_1 _13996_ (.A(_08893_),
    .X(_00155_));
 sky130_fd_sc_hd__buf_6 _13997_ (.A(_08547_),
    .X(_08894_));
 sky130_fd_sc_hd__mux2_1 _13998_ (.A0(_08894_),
    .A1(\cur_mb_mem[0][5] ),
    .S(_08884_),
    .X(_08895_));
 sky130_fd_sc_hd__clkbuf_1 _13999_ (.A(_08895_),
    .X(_00156_));
 sky130_fd_sc_hd__clkbuf_8 _14000_ (.A(_08550_),
    .X(_08896_));
 sky130_fd_sc_hd__mux2_1 _14001_ (.A0(_08896_),
    .A1(net1818),
    .S(_08884_),
    .X(_08897_));
 sky130_fd_sc_hd__clkbuf_1 _14002_ (.A(_08897_),
    .X(_00157_));
 sky130_fd_sc_hd__clkbuf_8 _14003_ (.A(_08553_),
    .X(_08898_));
 sky130_fd_sc_hd__mux2_1 _14004_ (.A0(_08898_),
    .A1(\cur_mb_mem[0][7] ),
    .S(_08884_),
    .X(_08899_));
 sky130_fd_sc_hd__clkbuf_1 _14005_ (.A(_08899_),
    .X(_00158_));
 sky130_fd_sc_hd__buf_4 _14006_ (.A(_08880_),
    .X(_08900_));
 sky130_fd_sc_hd__buf_12 _14007_ (.A(_08900_),
    .X(_08901_));
 sky130_fd_sc_hd__buf_12 _14008_ (.A(_08901_),
    .X(_08902_));
 sky130_fd_sc_hd__nand2_8 _14009_ (.A(_05990_),
    .B(_08902_),
    .Y(_08903_));
 sky130_fd_sc_hd__mux2_1 _14010_ (.A0(_08879_),
    .A1(\cur_mb_mem[1][0] ),
    .S(_08903_),
    .X(_08904_));
 sky130_fd_sc_hd__clkbuf_1 _14011_ (.A(_08904_),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _14012_ (.A0(_08886_),
    .A1(\cur_mb_mem[1][1] ),
    .S(_08903_),
    .X(_08905_));
 sky130_fd_sc_hd__clkbuf_1 _14013_ (.A(_08905_),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _14014_ (.A0(_08888_),
    .A1(\cur_mb_mem[1][2] ),
    .S(_08903_),
    .X(_08906_));
 sky130_fd_sc_hd__clkbuf_1 _14015_ (.A(_08906_),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _14016_ (.A0(_08890_),
    .A1(net670),
    .S(_08903_),
    .X(_08907_));
 sky130_fd_sc_hd__clkbuf_1 _14017_ (.A(_08907_),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _14018_ (.A0(_08892_),
    .A1(net1655),
    .S(_08903_),
    .X(_08908_));
 sky130_fd_sc_hd__clkbuf_1 _14019_ (.A(_08908_),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _14020_ (.A0(_08894_),
    .A1(net1475),
    .S(_08903_),
    .X(_08909_));
 sky130_fd_sc_hd__clkbuf_1 _14021_ (.A(_08909_),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _14022_ (.A0(_08896_),
    .A1(net1721),
    .S(_08903_),
    .X(_08910_));
 sky130_fd_sc_hd__clkbuf_1 _14023_ (.A(_08910_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _14024_ (.A0(_08898_),
    .A1(\cur_mb_mem[1][7] ),
    .S(_08903_),
    .X(_08911_));
 sky130_fd_sc_hd__clkbuf_1 _14025_ (.A(_08911_),
    .X(_00166_));
 sky130_fd_sc_hd__or3_2 _14026_ (.A(_05899_),
    .B(_06265_),
    .C(_08532_),
    .X(_08912_));
 sky130_fd_sc_hd__buf_6 _14027_ (.A(_08912_),
    .X(_08913_));
 sky130_fd_sc_hd__mux2_1 _14028_ (.A0(_08879_),
    .A1(net1343),
    .S(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__clkbuf_1 _14029_ (.A(_08914_),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _14030_ (.A0(_08886_),
    .A1(net1701),
    .S(_08913_),
    .X(_08915_));
 sky130_fd_sc_hd__clkbuf_1 _14031_ (.A(_08915_),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _14032_ (.A0(_08888_),
    .A1(net1578),
    .S(_08913_),
    .X(_08916_));
 sky130_fd_sc_hd__clkbuf_1 _14033_ (.A(_08916_),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _14034_ (.A0(_08890_),
    .A1(net881),
    .S(_08913_),
    .X(_08917_));
 sky130_fd_sc_hd__clkbuf_1 _14035_ (.A(_08917_),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _14036_ (.A0(_08892_),
    .A1(net1588),
    .S(_08913_),
    .X(_08918_));
 sky130_fd_sc_hd__clkbuf_1 _14037_ (.A(_08918_),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _14038_ (.A0(_08894_),
    .A1(net1576),
    .S(_08913_),
    .X(_08919_));
 sky130_fd_sc_hd__clkbuf_1 _14039_ (.A(_08919_),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _14040_ (.A0(_08896_),
    .A1(net1545),
    .S(_08913_),
    .X(_08920_));
 sky130_fd_sc_hd__clkbuf_1 _14041_ (.A(_08920_),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _14042_ (.A0(_08898_),
    .A1(\cur_mb_mem[2][7] ),
    .S(_08913_),
    .X(_08921_));
 sky130_fd_sc_hd__clkbuf_1 _14043_ (.A(_08921_),
    .X(_00174_));
 sky130_fd_sc_hd__nand2_8 _14044_ (.A(_06290_),
    .B(_08902_),
    .Y(_08922_));
 sky130_fd_sc_hd__mux2_1 _14045_ (.A0(_08879_),
    .A1(net676),
    .S(_08922_),
    .X(_08923_));
 sky130_fd_sc_hd__clkbuf_1 _14046_ (.A(_08923_),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _14047_ (.A0(_08886_),
    .A1(net1551),
    .S(_08922_),
    .X(_08924_));
 sky130_fd_sc_hd__clkbuf_1 _14048_ (.A(_08924_),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _14049_ (.A0(_08888_),
    .A1(net1400),
    .S(_08922_),
    .X(_08925_));
 sky130_fd_sc_hd__clkbuf_1 _14050_ (.A(_08925_),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _14051_ (.A0(_08890_),
    .A1(net908),
    .S(_08922_),
    .X(_08926_));
 sky130_fd_sc_hd__clkbuf_1 _14052_ (.A(_08926_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _14053_ (.A0(_08892_),
    .A1(net1208),
    .S(_08922_),
    .X(_08927_));
 sky130_fd_sc_hd__clkbuf_1 _14054_ (.A(_08927_),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _14055_ (.A0(_08894_),
    .A1(net969),
    .S(_08922_),
    .X(_08928_));
 sky130_fd_sc_hd__clkbuf_1 _14056_ (.A(_08928_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _14057_ (.A0(_08896_),
    .A1(net1373),
    .S(_08922_),
    .X(_08929_));
 sky130_fd_sc_hd__clkbuf_1 _14058_ (.A(_08929_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _14059_ (.A0(_08898_),
    .A1(\cur_mb_mem[3][7] ),
    .S(_08922_),
    .X(_08930_));
 sky130_fd_sc_hd__clkbuf_1 _14060_ (.A(_08930_),
    .X(_00182_));
 sky130_fd_sc_hd__nand2_8 _14061_ (.A(_06162_),
    .B(_08902_),
    .Y(_08931_));
 sky130_fd_sc_hd__mux2_1 _14062_ (.A0(_08879_),
    .A1(net1404),
    .S(_08931_),
    .X(_08932_));
 sky130_fd_sc_hd__clkbuf_1 _14063_ (.A(_08932_),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _14064_ (.A0(_08886_),
    .A1(net1663),
    .S(_08931_),
    .X(_08933_));
 sky130_fd_sc_hd__clkbuf_1 _14065_ (.A(_08933_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _14066_ (.A0(_08888_),
    .A1(\cur_mb_mem[4][2] ),
    .S(_08931_),
    .X(_08934_));
 sky130_fd_sc_hd__clkbuf_1 _14067_ (.A(_08934_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _14068_ (.A0(_08890_),
    .A1(net1980),
    .S(_08931_),
    .X(_08935_));
 sky130_fd_sc_hd__clkbuf_1 _14069_ (.A(_08935_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _14070_ (.A0(_08892_),
    .A1(net1349),
    .S(_08931_),
    .X(_08936_));
 sky130_fd_sc_hd__clkbuf_1 _14071_ (.A(_08936_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _14072_ (.A0(_08894_),
    .A1(net1662),
    .S(_08931_),
    .X(_08937_));
 sky130_fd_sc_hd__clkbuf_1 _14073_ (.A(_08937_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _14074_ (.A0(_08896_),
    .A1(\cur_mb_mem[4][6] ),
    .S(_08931_),
    .X(_08938_));
 sky130_fd_sc_hd__clkbuf_1 _14075_ (.A(_08938_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _14076_ (.A0(_08898_),
    .A1(\cur_mb_mem[4][7] ),
    .S(_08931_),
    .X(_08939_));
 sky130_fd_sc_hd__clkbuf_1 _14077_ (.A(_08939_),
    .X(_00190_));
 sky130_fd_sc_hd__nand2_8 _14078_ (.A(_06157_),
    .B(_08902_),
    .Y(_08940_));
 sky130_fd_sc_hd__mux2_1 _14079_ (.A0(_08879_),
    .A1(net1754),
    .S(_08940_),
    .X(_08941_));
 sky130_fd_sc_hd__clkbuf_1 _14080_ (.A(_08941_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _14081_ (.A0(_08886_),
    .A1(net1978),
    .S(_08940_),
    .X(_08942_));
 sky130_fd_sc_hd__clkbuf_1 _14082_ (.A(_08942_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _14083_ (.A0(_08888_),
    .A1(net1780),
    .S(_08940_),
    .X(_08943_));
 sky130_fd_sc_hd__clkbuf_1 _14084_ (.A(_08943_),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _14085_ (.A0(_08890_),
    .A1(net1794),
    .S(_08940_),
    .X(_08944_));
 sky130_fd_sc_hd__clkbuf_1 _14086_ (.A(_08944_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _14087_ (.A0(_08892_),
    .A1(net529),
    .S(_08940_),
    .X(_08945_));
 sky130_fd_sc_hd__clkbuf_1 _14088_ (.A(_08945_),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _14089_ (.A0(_08894_),
    .A1(net734),
    .S(_08940_),
    .X(_08946_));
 sky130_fd_sc_hd__clkbuf_1 _14090_ (.A(_08946_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _14091_ (.A0(_08896_),
    .A1(net1304),
    .S(_08940_),
    .X(_08947_));
 sky130_fd_sc_hd__clkbuf_1 _14092_ (.A(_08947_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _14093_ (.A0(_08898_),
    .A1(net1234),
    .S(_08940_),
    .X(_08948_));
 sky130_fd_sc_hd__clkbuf_1 _14094_ (.A(_08948_),
    .X(_00198_));
 sky130_fd_sc_hd__nand2_8 _14095_ (.A(_06203_),
    .B(_08902_),
    .Y(_08949_));
 sky130_fd_sc_hd__mux2_1 _14096_ (.A0(_08879_),
    .A1(net1480),
    .S(_08949_),
    .X(_08950_));
 sky130_fd_sc_hd__clkbuf_1 _14097_ (.A(_08950_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _14098_ (.A0(_08886_),
    .A1(net1007),
    .S(_08949_),
    .X(_08951_));
 sky130_fd_sc_hd__clkbuf_1 _14099_ (.A(_08951_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _14100_ (.A0(_08888_),
    .A1(net1061),
    .S(_08949_),
    .X(_08952_));
 sky130_fd_sc_hd__clkbuf_1 _14101_ (.A(_08952_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _14102_ (.A0(_08890_),
    .A1(net1524),
    .S(_08949_),
    .X(_08953_));
 sky130_fd_sc_hd__clkbuf_1 _14103_ (.A(_08953_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _14104_ (.A0(_08892_),
    .A1(net728),
    .S(_08949_),
    .X(_08954_));
 sky130_fd_sc_hd__clkbuf_1 _14105_ (.A(_08954_),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _14106_ (.A0(_08894_),
    .A1(net1027),
    .S(_08949_),
    .X(_08955_));
 sky130_fd_sc_hd__clkbuf_1 _14107_ (.A(_08955_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _14108_ (.A0(_08896_),
    .A1(net1363),
    .S(_08949_),
    .X(_08956_));
 sky130_fd_sc_hd__clkbuf_1 _14109_ (.A(_08956_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _14110_ (.A0(_08898_),
    .A1(net1348),
    .S(_08949_),
    .X(_08957_));
 sky130_fd_sc_hd__clkbuf_1 _14111_ (.A(_08957_),
    .X(_00206_));
 sky130_fd_sc_hd__buf_6 _14112_ (.A(_08900_),
    .X(_08958_));
 sky130_fd_sc_hd__and3_1 _14113_ (.A(_06113_),
    .B(_08839_),
    .C(_08958_),
    .X(_08959_));
 sky130_fd_sc_hd__buf_6 _14114_ (.A(_08959_),
    .X(_08960_));
 sky130_fd_sc_hd__mux2_1 _14115_ (.A0(net358),
    .A1(_08531_),
    .S(_08960_),
    .X(_08961_));
 sky130_fd_sc_hd__clkbuf_1 _14116_ (.A(_08961_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _14117_ (.A0(net506),
    .A1(_08536_),
    .S(_08960_),
    .X(_08962_));
 sky130_fd_sc_hd__clkbuf_1 _14118_ (.A(_08962_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _14119_ (.A0(net390),
    .A1(_08539_),
    .S(_08960_),
    .X(_08963_));
 sky130_fd_sc_hd__clkbuf_1 _14120_ (.A(_08963_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _14121_ (.A0(net453),
    .A1(_08542_),
    .S(_08960_),
    .X(_08964_));
 sky130_fd_sc_hd__clkbuf_1 _14122_ (.A(_08964_),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _14123_ (.A0(net410),
    .A1(_08545_),
    .S(_08960_),
    .X(_08965_));
 sky130_fd_sc_hd__clkbuf_1 _14124_ (.A(_08965_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _14125_ (.A0(net368),
    .A1(_08548_),
    .S(_08960_),
    .X(_08966_));
 sky130_fd_sc_hd__clkbuf_1 _14126_ (.A(_08966_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _14127_ (.A0(net1255),
    .A1(_08551_),
    .S(_08960_),
    .X(_08967_));
 sky130_fd_sc_hd__clkbuf_1 _14128_ (.A(_08967_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _14129_ (.A0(net1565),
    .A1(_08554_),
    .S(_08960_),
    .X(_08968_));
 sky130_fd_sc_hd__clkbuf_1 _14130_ (.A(_08968_),
    .X(_00214_));
 sky130_fd_sc_hd__nand2_8 _14131_ (.A(_06277_),
    .B(_08902_),
    .Y(_08969_));
 sky130_fd_sc_hd__mux2_1 _14132_ (.A0(_08879_),
    .A1(net1311),
    .S(_08969_),
    .X(_08970_));
 sky130_fd_sc_hd__clkbuf_1 _14133_ (.A(_08970_),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _14134_ (.A0(_08886_),
    .A1(net1134),
    .S(_08969_),
    .X(_08971_));
 sky130_fd_sc_hd__clkbuf_1 _14135_ (.A(_08971_),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _14136_ (.A0(_08888_),
    .A1(net1376),
    .S(_08969_),
    .X(_08972_));
 sky130_fd_sc_hd__clkbuf_1 _14137_ (.A(_08972_),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _14138_ (.A0(_08890_),
    .A1(net1036),
    .S(_08969_),
    .X(_08973_));
 sky130_fd_sc_hd__clkbuf_1 _14139_ (.A(_08973_),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _14140_ (.A0(_08892_),
    .A1(net912),
    .S(_08969_),
    .X(_08974_));
 sky130_fd_sc_hd__clkbuf_1 _14141_ (.A(_08974_),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _14142_ (.A0(_08894_),
    .A1(net1160),
    .S(_08969_),
    .X(_08975_));
 sky130_fd_sc_hd__clkbuf_1 _14143_ (.A(_08975_),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _14144_ (.A0(_08896_),
    .A1(net1405),
    .S(_08969_),
    .X(_08976_));
 sky130_fd_sc_hd__clkbuf_1 _14145_ (.A(_08976_),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _14146_ (.A0(_08898_),
    .A1(net887),
    .S(_08969_),
    .X(_08977_));
 sky130_fd_sc_hd__clkbuf_1 _14147_ (.A(_08977_),
    .X(_00222_));
 sky130_fd_sc_hd__buf_8 _14148_ (.A(_05912_),
    .X(_08978_));
 sky130_fd_sc_hd__buf_12 _14149_ (.A(_08958_),
    .X(_08979_));
 sky130_fd_sc_hd__nand3_4 _14150_ (.A(_06113_),
    .B(_08978_),
    .C(_08979_),
    .Y(_08980_));
 sky130_fd_sc_hd__mux2_1 _14151_ (.A0(_08879_),
    .A1(net860),
    .S(net216),
    .X(_08981_));
 sky130_fd_sc_hd__clkbuf_1 _14152_ (.A(_08981_),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _14153_ (.A0(_08886_),
    .A1(net716),
    .S(net216),
    .X(_08982_));
 sky130_fd_sc_hd__clkbuf_1 _14154_ (.A(_08982_),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _14155_ (.A0(_08888_),
    .A1(net1260),
    .S(net216),
    .X(_08983_));
 sky130_fd_sc_hd__clkbuf_1 _14156_ (.A(_08983_),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _14157_ (.A0(_08890_),
    .A1(net915),
    .S(net216),
    .X(_08984_));
 sky130_fd_sc_hd__clkbuf_1 _14158_ (.A(_08984_),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _14159_ (.A0(_08892_),
    .A1(net694),
    .S(_08980_),
    .X(_08985_));
 sky130_fd_sc_hd__clkbuf_1 _14160_ (.A(_08985_),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _14161_ (.A0(_08894_),
    .A1(net1079),
    .S(_08980_),
    .X(_08986_));
 sky130_fd_sc_hd__clkbuf_1 _14162_ (.A(_08986_),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _14163_ (.A0(_08896_),
    .A1(net449),
    .S(net216),
    .X(_08987_));
 sky130_fd_sc_hd__clkbuf_1 _14164_ (.A(_08987_),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _14165_ (.A0(_08898_),
    .A1(net888),
    .S(net216),
    .X(_08988_));
 sky130_fd_sc_hd__clkbuf_1 _14166_ (.A(_08988_),
    .X(_00230_));
 sky130_fd_sc_hd__nand2_8 _14167_ (.A(_06408_),
    .B(_08902_),
    .Y(_08989_));
 sky130_fd_sc_hd__mux2_1 _14168_ (.A0(_08879_),
    .A1(net1439),
    .S(_08989_),
    .X(_08990_));
 sky130_fd_sc_hd__clkbuf_1 _14169_ (.A(_08990_),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _14170_ (.A0(_08886_),
    .A1(net1503),
    .S(_08989_),
    .X(_08991_));
 sky130_fd_sc_hd__clkbuf_1 _14171_ (.A(_08991_),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _14172_ (.A0(_08888_),
    .A1(net1226),
    .S(_08989_),
    .X(_08992_));
 sky130_fd_sc_hd__clkbuf_1 _14173_ (.A(_08992_),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _14174_ (.A0(_08890_),
    .A1(net1802),
    .S(_08989_),
    .X(_08993_));
 sky130_fd_sc_hd__clkbuf_1 _14175_ (.A(_08993_),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _14176_ (.A0(_08892_),
    .A1(net1431),
    .S(_08989_),
    .X(_08994_));
 sky130_fd_sc_hd__clkbuf_1 _14177_ (.A(_08994_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _14178_ (.A0(_08894_),
    .A1(net1497),
    .S(_08989_),
    .X(_08995_));
 sky130_fd_sc_hd__clkbuf_1 _14179_ (.A(_08995_),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _14180_ (.A0(_08896_),
    .A1(net1198),
    .S(_08989_),
    .X(_08996_));
 sky130_fd_sc_hd__clkbuf_1 _14181_ (.A(_08996_),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _14182_ (.A0(_08898_),
    .A1(net1359),
    .S(_08989_),
    .X(_08997_));
 sky130_fd_sc_hd__clkbuf_1 _14183_ (.A(_08997_),
    .X(_00238_));
 sky130_fd_sc_hd__and3_1 _14184_ (.A(_06113_),
    .B(_06049_),
    .C(_08958_),
    .X(_08998_));
 sky130_fd_sc_hd__buf_4 _14185_ (.A(_08998_),
    .X(_08999_));
 sky130_fd_sc_hd__mux2_1 _14186_ (.A0(net925),
    .A1(_08531_),
    .S(_08999_),
    .X(_09000_));
 sky130_fd_sc_hd__clkbuf_1 _14187_ (.A(_09000_),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _14188_ (.A0(net1838),
    .A1(_08536_),
    .S(_08999_),
    .X(_09001_));
 sky130_fd_sc_hd__clkbuf_1 _14189_ (.A(_09001_),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _14190_ (.A0(net1396),
    .A1(_08539_),
    .S(_08999_),
    .X(_09002_));
 sky130_fd_sc_hd__clkbuf_1 _14191_ (.A(_09002_),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _14192_ (.A0(net1370),
    .A1(_08542_),
    .S(_08999_),
    .X(_09003_));
 sky130_fd_sc_hd__clkbuf_1 _14193_ (.A(_09003_),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _14194_ (.A0(net1446),
    .A1(_08545_),
    .S(_08999_),
    .X(_09004_));
 sky130_fd_sc_hd__clkbuf_1 _14195_ (.A(_09004_),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _14196_ (.A0(net1291),
    .A1(_08548_),
    .S(_08999_),
    .X(_09005_));
 sky130_fd_sc_hd__clkbuf_1 _14197_ (.A(_09005_),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _14198_ (.A0(net1777),
    .A1(_08551_),
    .S(_08999_),
    .X(_09006_));
 sky130_fd_sc_hd__clkbuf_1 _14199_ (.A(_09006_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _14200_ (.A0(net839),
    .A1(_08554_),
    .S(_08999_),
    .X(_09007_));
 sky130_fd_sc_hd__clkbuf_1 _14201_ (.A(_09007_),
    .X(_00246_));
 sky130_fd_sc_hd__clkbuf_16 _14202_ (.A(_08530_),
    .X(_09008_));
 sky130_fd_sc_hd__nand2_8 _14203_ (.A(_05928_),
    .B(_08902_),
    .Y(_09009_));
 sky130_fd_sc_hd__mux2_1 _14204_ (.A0(_09008_),
    .A1(net1623),
    .S(_09009_),
    .X(_09010_));
 sky130_fd_sc_hd__clkbuf_1 _14205_ (.A(_09010_),
    .X(_00247_));
 sky130_fd_sc_hd__buf_6 _14206_ (.A(_08535_),
    .X(_09011_));
 sky130_fd_sc_hd__mux2_1 _14207_ (.A0(_09011_),
    .A1(net1202),
    .S(_09009_),
    .X(_09012_));
 sky130_fd_sc_hd__clkbuf_1 _14208_ (.A(_09012_),
    .X(_00248_));
 sky130_fd_sc_hd__clkbuf_16 _14209_ (.A(_08538_),
    .X(_09013_));
 sky130_fd_sc_hd__mux2_1 _14210_ (.A0(_09013_),
    .A1(net1854),
    .S(_09009_),
    .X(_09014_));
 sky130_fd_sc_hd__clkbuf_1 _14211_ (.A(_09014_),
    .X(_00249_));
 sky130_fd_sc_hd__clkbuf_16 _14212_ (.A(_08541_),
    .X(_09015_));
 sky130_fd_sc_hd__mux2_1 _14213_ (.A0(_09015_),
    .A1(net1720),
    .S(_09009_),
    .X(_09016_));
 sky130_fd_sc_hd__clkbuf_1 _14214_ (.A(_09016_),
    .X(_00250_));
 sky130_fd_sc_hd__buf_6 _14215_ (.A(_08544_),
    .X(_09017_));
 sky130_fd_sc_hd__mux2_1 _14216_ (.A0(_09017_),
    .A1(net1244),
    .S(_09009_),
    .X(_09018_));
 sky130_fd_sc_hd__clkbuf_1 _14217_ (.A(_09018_),
    .X(_00251_));
 sky130_fd_sc_hd__buf_6 _14218_ (.A(_08547_),
    .X(_09019_));
 sky130_fd_sc_hd__mux2_1 _14219_ (.A0(_09019_),
    .A1(net1212),
    .S(_09009_),
    .X(_09020_));
 sky130_fd_sc_hd__clkbuf_1 _14220_ (.A(_09020_),
    .X(_00252_));
 sky130_fd_sc_hd__clkbuf_8 _14221_ (.A(_08550_),
    .X(_09021_));
 sky130_fd_sc_hd__mux2_1 _14222_ (.A0(_09021_),
    .A1(\cur_mb_mem[12][6] ),
    .S(_09009_),
    .X(_09022_));
 sky130_fd_sc_hd__clkbuf_1 _14223_ (.A(_09022_),
    .X(_00253_));
 sky130_fd_sc_hd__buf_6 _14224_ (.A(_08553_),
    .X(_09023_));
 sky130_fd_sc_hd__mux2_1 _14225_ (.A0(_09023_),
    .A1(net1152),
    .S(_09009_),
    .X(_09024_));
 sky130_fd_sc_hd__clkbuf_1 _14226_ (.A(_09024_),
    .X(_00254_));
 sky130_fd_sc_hd__buf_6 _14227_ (.A(_05961_),
    .X(_09025_));
 sky130_fd_sc_hd__and3_1 _14228_ (.A(_06113_),
    .B(_09025_),
    .C(_08958_),
    .X(_09026_));
 sky130_fd_sc_hd__buf_4 _14229_ (.A(_09026_),
    .X(_09027_));
 sky130_fd_sc_hd__mux2_1 _14230_ (.A0(net1930),
    .A1(_08531_),
    .S(_09027_),
    .X(_09028_));
 sky130_fd_sc_hd__clkbuf_1 _14231_ (.A(_09028_),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _14232_ (.A0(net597),
    .A1(_08536_),
    .S(_09027_),
    .X(_09029_));
 sky130_fd_sc_hd__clkbuf_1 _14233_ (.A(_09029_),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _14234_ (.A0(net1730),
    .A1(_08539_),
    .S(_09027_),
    .X(_09030_));
 sky130_fd_sc_hd__clkbuf_1 _14235_ (.A(_09030_),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _14236_ (.A0(net1899),
    .A1(_08542_),
    .S(_09027_),
    .X(_09031_));
 sky130_fd_sc_hd__clkbuf_1 _14237_ (.A(_09031_),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _14238_ (.A0(net1355),
    .A1(_08545_),
    .S(_09027_),
    .X(_09032_));
 sky130_fd_sc_hd__clkbuf_1 _14239_ (.A(_09032_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _14240_ (.A0(net1215),
    .A1(_08548_),
    .S(_09027_),
    .X(_09033_));
 sky130_fd_sc_hd__clkbuf_1 _14241_ (.A(_09033_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _14242_ (.A0(net740),
    .A1(_08551_),
    .S(_09027_),
    .X(_09034_));
 sky130_fd_sc_hd__clkbuf_1 _14243_ (.A(_09034_),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _14244_ (.A0(net639),
    .A1(_08554_),
    .S(_09027_),
    .X(_09035_));
 sky130_fd_sc_hd__clkbuf_1 _14245_ (.A(_09035_),
    .X(_00262_));
 sky130_fd_sc_hd__buf_6 _14246_ (.A(_06025_),
    .X(_09036_));
 sky130_fd_sc_hd__clkbuf_2 _14247_ (.A(_08900_),
    .X(_09037_));
 sky130_fd_sc_hd__and3_1 _14248_ (.A(_06113_),
    .B(_09036_),
    .C(_09037_),
    .X(_09038_));
 sky130_fd_sc_hd__buf_8 _14249_ (.A(_09038_),
    .X(_09039_));
 sky130_fd_sc_hd__mux2_1 _14250_ (.A0(net1142),
    .A1(_08531_),
    .S(_09039_),
    .X(_09040_));
 sky130_fd_sc_hd__clkbuf_1 _14251_ (.A(_09040_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _14252_ (.A0(net800),
    .A1(_08536_),
    .S(_09039_),
    .X(_09041_));
 sky130_fd_sc_hd__clkbuf_1 _14253_ (.A(_09041_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _14254_ (.A0(net1689),
    .A1(_08539_),
    .S(_09039_),
    .X(_09042_));
 sky130_fd_sc_hd__clkbuf_1 _14255_ (.A(_09042_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _14256_ (.A0(net935),
    .A1(_08542_),
    .S(_09039_),
    .X(_09043_));
 sky130_fd_sc_hd__clkbuf_1 _14257_ (.A(_09043_),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _14258_ (.A0(net1337),
    .A1(_08545_),
    .S(_09039_),
    .X(_09044_));
 sky130_fd_sc_hd__clkbuf_1 _14259_ (.A(_09044_),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _14260_ (.A0(net1043),
    .A1(_08548_),
    .S(_09039_),
    .X(_09045_));
 sky130_fd_sc_hd__clkbuf_1 _14261_ (.A(_09045_),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _14262_ (.A0(net754),
    .A1(_08551_),
    .S(_09039_),
    .X(_09046_));
 sky130_fd_sc_hd__clkbuf_1 _14263_ (.A(_09046_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _14264_ (.A0(net1016),
    .A1(_08554_),
    .S(_09039_),
    .X(_09047_));
 sky130_fd_sc_hd__clkbuf_1 _14265_ (.A(_09047_),
    .X(_00270_));
 sky130_fd_sc_hd__nand2_8 _14266_ (.A(_06295_),
    .B(_08902_),
    .Y(_09048_));
 sky130_fd_sc_hd__mux2_1 _14267_ (.A0(_09008_),
    .A1(net897),
    .S(_09048_),
    .X(_09049_));
 sky130_fd_sc_hd__clkbuf_1 _14268_ (.A(_09049_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _14269_ (.A0(_09011_),
    .A1(net1305),
    .S(_09048_),
    .X(_09050_));
 sky130_fd_sc_hd__clkbuf_1 _14270_ (.A(_09050_),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _14271_ (.A0(_09013_),
    .A1(net1335),
    .S(_09048_),
    .X(_09051_));
 sky130_fd_sc_hd__clkbuf_1 _14272_ (.A(_09051_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _14273_ (.A0(_09015_),
    .A1(net868),
    .S(_09048_),
    .X(_09052_));
 sky130_fd_sc_hd__clkbuf_1 _14274_ (.A(_09052_),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _14275_ (.A0(_09017_),
    .A1(\cur_mb_mem[15][4] ),
    .S(_09048_),
    .X(_09053_));
 sky130_fd_sc_hd__clkbuf_1 _14276_ (.A(_09053_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _14277_ (.A0(_09019_),
    .A1(\cur_mb_mem[15][5] ),
    .S(_09048_),
    .X(_09054_));
 sky130_fd_sc_hd__clkbuf_1 _14278_ (.A(_09054_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _14279_ (.A0(_09021_),
    .A1(net1085),
    .S(_09048_),
    .X(_09055_));
 sky130_fd_sc_hd__clkbuf_1 _14280_ (.A(_09055_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _14281_ (.A0(_09023_),
    .A1(net1426),
    .S(_09048_),
    .X(_09056_));
 sky130_fd_sc_hd__clkbuf_1 _14282_ (.A(_09056_),
    .X(_00278_));
 sky130_fd_sc_hd__nand2_8 _14283_ (.A(_05976_),
    .B(_08883_),
    .Y(_09057_));
 sky130_fd_sc_hd__mux2_1 _14284_ (.A0(_09008_),
    .A1(net739),
    .S(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__clkbuf_1 _14285_ (.A(_09058_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _14286_ (.A0(_09011_),
    .A1(net620),
    .S(_09057_),
    .X(_09059_));
 sky130_fd_sc_hd__clkbuf_1 _14287_ (.A(_09059_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _14288_ (.A0(_09013_),
    .A1(net1393),
    .S(_09057_),
    .X(_09060_));
 sky130_fd_sc_hd__clkbuf_1 _14289_ (.A(_09060_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _14290_ (.A0(_09015_),
    .A1(net579),
    .S(_09057_),
    .X(_09061_));
 sky130_fd_sc_hd__clkbuf_1 _14291_ (.A(_09061_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _14292_ (.A0(_09017_),
    .A1(net810),
    .S(_09057_),
    .X(_09062_));
 sky130_fd_sc_hd__clkbuf_1 _14293_ (.A(_09062_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _14294_ (.A0(_09019_),
    .A1(net674),
    .S(_09057_),
    .X(_09063_));
 sky130_fd_sc_hd__clkbuf_1 _14295_ (.A(_09063_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _14296_ (.A0(_09021_),
    .A1(net1166),
    .S(_09057_),
    .X(_09064_));
 sky130_fd_sc_hd__clkbuf_1 _14297_ (.A(_09064_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _14298_ (.A0(_09023_),
    .A1(net1530),
    .S(_09057_),
    .X(_09065_));
 sky130_fd_sc_hd__clkbuf_1 _14299_ (.A(_09065_),
    .X(_00286_));
 sky130_fd_sc_hd__nand2_8 _14300_ (.A(_06318_),
    .B(_08902_),
    .Y(_09066_));
 sky130_fd_sc_hd__mux2_1 _14301_ (.A0(_09008_),
    .A1(net686),
    .S(_09066_),
    .X(_09067_));
 sky130_fd_sc_hd__clkbuf_1 _14302_ (.A(_09067_),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _14303_ (.A0(_09011_),
    .A1(net657),
    .S(_09066_),
    .X(_09068_));
 sky130_fd_sc_hd__clkbuf_1 _14304_ (.A(_09068_),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _14305_ (.A0(_09013_),
    .A1(net792),
    .S(_09066_),
    .X(_09069_));
 sky130_fd_sc_hd__clkbuf_1 _14306_ (.A(_09069_),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _14307_ (.A0(_09015_),
    .A1(net1394),
    .S(_09066_),
    .X(_09070_));
 sky130_fd_sc_hd__clkbuf_1 _14308_ (.A(_09070_),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _14309_ (.A0(_09017_),
    .A1(net1424),
    .S(_09066_),
    .X(_09071_));
 sky130_fd_sc_hd__clkbuf_1 _14310_ (.A(_09071_),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _14311_ (.A0(_09019_),
    .A1(net1476),
    .S(_09066_),
    .X(_09072_));
 sky130_fd_sc_hd__clkbuf_1 _14312_ (.A(_09072_),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _14313_ (.A0(_09021_),
    .A1(\cur_mb_mem[17][6] ),
    .S(_09066_),
    .X(_09073_));
 sky130_fd_sc_hd__clkbuf_1 _14314_ (.A(_09073_),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _14315_ (.A0(_09023_),
    .A1(net1412),
    .S(_09066_),
    .X(_09074_));
 sky130_fd_sc_hd__clkbuf_1 _14316_ (.A(_09074_),
    .X(_00294_));
 sky130_fd_sc_hd__or3_1 _14317_ (.A(_06265_),
    .B(_06177_),
    .C(_08532_),
    .X(_09075_));
 sky130_fd_sc_hd__buf_8 _14318_ (.A(_09075_),
    .X(_09076_));
 sky130_fd_sc_hd__mux2_1 _14319_ (.A0(_09008_),
    .A1(net1227),
    .S(_09076_),
    .X(_09077_));
 sky130_fd_sc_hd__clkbuf_1 _14320_ (.A(_09077_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _14321_ (.A0(_09011_),
    .A1(net614),
    .S(_09076_),
    .X(_09078_));
 sky130_fd_sc_hd__clkbuf_1 _14322_ (.A(_09078_),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _14323_ (.A0(_09013_),
    .A1(net932),
    .S(_09076_),
    .X(_09079_));
 sky130_fd_sc_hd__clkbuf_1 _14324_ (.A(_09079_),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _14325_ (.A0(_09015_),
    .A1(\cur_mb_mem[18][3] ),
    .S(_09076_),
    .X(_09080_));
 sky130_fd_sc_hd__clkbuf_1 _14326_ (.A(_09080_),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _14327_ (.A0(_09017_),
    .A1(net822),
    .S(_09076_),
    .X(_09081_));
 sky130_fd_sc_hd__clkbuf_1 _14328_ (.A(_09081_),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _14329_ (.A0(_09019_),
    .A1(net628),
    .S(_09076_),
    .X(_09082_));
 sky130_fd_sc_hd__clkbuf_1 _14330_ (.A(_09082_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _14331_ (.A0(_09021_),
    .A1(net1124),
    .S(_09076_),
    .X(_09083_));
 sky130_fd_sc_hd__clkbuf_1 _14332_ (.A(_09083_),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _14333_ (.A0(_09023_),
    .A1(net1267),
    .S(_09076_),
    .X(_09084_));
 sky130_fd_sc_hd__clkbuf_1 _14334_ (.A(_09084_),
    .X(_00302_));
 sky130_fd_sc_hd__buf_12 _14335_ (.A(_08901_),
    .X(_09085_));
 sky130_fd_sc_hd__nand2_8 _14336_ (.A(_06282_),
    .B(_09085_),
    .Y(_09086_));
 sky130_fd_sc_hd__mux2_1 _14337_ (.A0(_09008_),
    .A1(net1379),
    .S(_09086_),
    .X(_09087_));
 sky130_fd_sc_hd__clkbuf_1 _14338_ (.A(_09087_),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _14339_ (.A0(_09011_),
    .A1(net1464),
    .S(_09086_),
    .X(_09088_));
 sky130_fd_sc_hd__clkbuf_1 _14340_ (.A(_09088_),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _14341_ (.A0(_09013_),
    .A1(net1278),
    .S(_09086_),
    .X(_09089_));
 sky130_fd_sc_hd__clkbuf_1 _14342_ (.A(_09089_),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _14343_ (.A0(_09015_),
    .A1(net1444),
    .S(_09086_),
    .X(_09090_));
 sky130_fd_sc_hd__clkbuf_1 _14344_ (.A(_09090_),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _14345_ (.A0(_09017_),
    .A1(net1187),
    .S(_09086_),
    .X(_09091_));
 sky130_fd_sc_hd__clkbuf_1 _14346_ (.A(_09091_),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _14347_ (.A0(_09019_),
    .A1(net1395),
    .S(_09086_),
    .X(_09092_));
 sky130_fd_sc_hd__clkbuf_1 _14348_ (.A(_09092_),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _14349_ (.A0(_09021_),
    .A1(net1163),
    .S(_09086_),
    .X(_09093_));
 sky130_fd_sc_hd__clkbuf_1 _14350_ (.A(_09093_),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _14351_ (.A0(_09023_),
    .A1(net1275),
    .S(_09086_),
    .X(_09094_));
 sky130_fd_sc_hd__clkbuf_1 _14352_ (.A(_09094_),
    .X(_00310_));
 sky130_fd_sc_hd__or3_1 _14353_ (.A(_06161_),
    .B(_06177_),
    .C(_08532_),
    .X(_09095_));
 sky130_fd_sc_hd__buf_4 _14354_ (.A(_09095_),
    .X(_09096_));
 sky130_fd_sc_hd__mux2_1 _14355_ (.A0(_09008_),
    .A1(net1171),
    .S(_09096_),
    .X(_09097_));
 sky130_fd_sc_hd__clkbuf_1 _14356_ (.A(_09097_),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _14357_ (.A0(_09011_),
    .A1(net801),
    .S(_09096_),
    .X(_09098_));
 sky130_fd_sc_hd__clkbuf_1 _14358_ (.A(_09098_),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _14359_ (.A0(_09013_),
    .A1(net1225),
    .S(_09096_),
    .X(_09099_));
 sky130_fd_sc_hd__clkbuf_1 _14360_ (.A(_09099_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _14361_ (.A0(_09015_),
    .A1(net1514),
    .S(_09096_),
    .X(_09100_));
 sky130_fd_sc_hd__clkbuf_1 _14362_ (.A(_09100_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _14363_ (.A0(_09017_),
    .A1(net1203),
    .S(_09096_),
    .X(_09101_));
 sky130_fd_sc_hd__clkbuf_1 _14364_ (.A(_09101_),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _14365_ (.A0(_09019_),
    .A1(net1483),
    .S(_09096_),
    .X(_09102_));
 sky130_fd_sc_hd__clkbuf_1 _14366_ (.A(_09102_),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _14367_ (.A0(_09021_),
    .A1(net1008),
    .S(_09096_),
    .X(_09103_));
 sky130_fd_sc_hd__clkbuf_1 _14368_ (.A(_09103_),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _14369_ (.A0(_09023_),
    .A1(net1591),
    .S(_09096_),
    .X(_09104_));
 sky130_fd_sc_hd__clkbuf_1 _14370_ (.A(_09104_),
    .X(_00318_));
 sky130_fd_sc_hd__nand2_8 _14371_ (.A(_06236_),
    .B(_09085_),
    .Y(_09105_));
 sky130_fd_sc_hd__mux2_1 _14372_ (.A0(_09008_),
    .A1(net862),
    .S(_09105_),
    .X(_09106_));
 sky130_fd_sc_hd__clkbuf_1 _14373_ (.A(_09106_),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _14374_ (.A0(_09011_),
    .A1(net1350),
    .S(_09105_),
    .X(_09107_));
 sky130_fd_sc_hd__clkbuf_1 _14375_ (.A(_09107_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _14376_ (.A0(_09013_),
    .A1(net720),
    .S(_09105_),
    .X(_09108_));
 sky130_fd_sc_hd__clkbuf_1 _14377_ (.A(_09108_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _14378_ (.A0(_09015_),
    .A1(net793),
    .S(_09105_),
    .X(_09109_));
 sky130_fd_sc_hd__clkbuf_1 _14379_ (.A(_09109_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _14380_ (.A0(_09017_),
    .A1(net1078),
    .S(_09105_),
    .X(_09110_));
 sky130_fd_sc_hd__clkbuf_1 _14381_ (.A(_09110_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _14382_ (.A0(_09019_),
    .A1(net1518),
    .S(_09105_),
    .X(_09111_));
 sky130_fd_sc_hd__clkbuf_1 _14383_ (.A(_09111_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _14384_ (.A0(_09021_),
    .A1(net1274),
    .S(_09105_),
    .X(_09112_));
 sky130_fd_sc_hd__clkbuf_1 _14385_ (.A(_09112_),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _14386_ (.A0(_09023_),
    .A1(net1101),
    .S(_09105_),
    .X(_09113_));
 sky130_fd_sc_hd__clkbuf_1 _14387_ (.A(_09113_),
    .X(_00326_));
 sky130_fd_sc_hd__nand2_8 _14388_ (.A(_06242_),
    .B(_09085_),
    .Y(_09114_));
 sky130_fd_sc_hd__mux2_1 _14389_ (.A0(_09008_),
    .A1(net1589),
    .S(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__clkbuf_1 _14390_ (.A(_09115_),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _14391_ (.A0(_09011_),
    .A1(net1290),
    .S(_09114_),
    .X(_09116_));
 sky130_fd_sc_hd__clkbuf_1 _14392_ (.A(_09116_),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _14393_ (.A0(_09013_),
    .A1(net1534),
    .S(_09114_),
    .X(_09117_));
 sky130_fd_sc_hd__clkbuf_1 _14394_ (.A(_09117_),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _14395_ (.A0(_09015_),
    .A1(net1493),
    .S(_09114_),
    .X(_09118_));
 sky130_fd_sc_hd__clkbuf_1 _14396_ (.A(_09118_),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _14397_ (.A0(_09017_),
    .A1(net831),
    .S(_09114_),
    .X(_09119_));
 sky130_fd_sc_hd__clkbuf_1 _14398_ (.A(_09119_),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _14399_ (.A0(_09019_),
    .A1(net930),
    .S(_09114_),
    .X(_09120_));
 sky130_fd_sc_hd__clkbuf_1 _14400_ (.A(_09120_),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _14401_ (.A0(_09021_),
    .A1(net1334),
    .S(_09114_),
    .X(_09121_));
 sky130_fd_sc_hd__clkbuf_1 _14402_ (.A(_09121_),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _14403_ (.A0(_09023_),
    .A1(net1246),
    .S(_09114_),
    .X(_09122_));
 sky130_fd_sc_hd__clkbuf_1 _14404_ (.A(_09122_),
    .X(_00334_));
 sky130_fd_sc_hd__nand3_4 _14405_ (.A(_08839_),
    .B(_05976_),
    .C(_08979_),
    .Y(_09123_));
 sky130_fd_sc_hd__mux2_1 _14406_ (.A0(_09008_),
    .A1(net591),
    .S(_09123_),
    .X(_09124_));
 sky130_fd_sc_hd__clkbuf_1 _14407_ (.A(_09124_),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _14408_ (.A0(_09011_),
    .A1(net838),
    .S(net215),
    .X(_09125_));
 sky130_fd_sc_hd__clkbuf_1 _14409_ (.A(_09125_),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _14410_ (.A0(_09013_),
    .A1(net913),
    .S(net215),
    .X(_09126_));
 sky130_fd_sc_hd__clkbuf_1 _14411_ (.A(_09126_),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _14412_ (.A0(_09015_),
    .A1(net779),
    .S(net215),
    .X(_09127_));
 sky130_fd_sc_hd__clkbuf_1 _14413_ (.A(_09127_),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _14414_ (.A0(_09017_),
    .A1(net1090),
    .S(net215),
    .X(_09128_));
 sky130_fd_sc_hd__clkbuf_1 _14415_ (.A(_09128_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _14416_ (.A0(_09019_),
    .A1(net997),
    .S(net215),
    .X(_09129_));
 sky130_fd_sc_hd__clkbuf_1 _14417_ (.A(_09129_),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _14418_ (.A0(_09021_),
    .A1(net1842),
    .S(_09123_),
    .X(_09130_));
 sky130_fd_sc_hd__clkbuf_1 _14419_ (.A(_09130_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _14420_ (.A0(_09023_),
    .A1(net1499),
    .S(_09123_),
    .X(_09131_));
 sky130_fd_sc_hd__clkbuf_1 _14421_ (.A(_09131_),
    .X(_00342_));
 sky130_fd_sc_hd__buf_8 _14422_ (.A(net97),
    .X(_09132_));
 sky130_fd_sc_hd__buf_4 _14423_ (.A(_09132_),
    .X(_09133_));
 sky130_fd_sc_hd__nand2_4 _14424_ (.A(_06285_),
    .B(_09085_),
    .Y(_09134_));
 sky130_fd_sc_hd__mux2_1 _14425_ (.A0(_09133_),
    .A1(net1603),
    .S(_09134_),
    .X(_09135_));
 sky130_fd_sc_hd__clkbuf_1 _14426_ (.A(_09135_),
    .X(_00343_));
 sky130_fd_sc_hd__buf_6 _14427_ (.A(net98),
    .X(_09136_));
 sky130_fd_sc_hd__buf_4 _14428_ (.A(_09136_),
    .X(_09137_));
 sky130_fd_sc_hd__mux2_1 _14429_ (.A0(_09137_),
    .A1(net1540),
    .S(_09134_),
    .X(_09138_));
 sky130_fd_sc_hd__clkbuf_1 _14430_ (.A(_09138_),
    .X(_00344_));
 sky130_fd_sc_hd__buf_6 _14431_ (.A(net99),
    .X(_09139_));
 sky130_fd_sc_hd__buf_4 _14432_ (.A(_09139_),
    .X(_09140_));
 sky130_fd_sc_hd__mux2_1 _14433_ (.A0(_09140_),
    .A1(net1738),
    .S(_09134_),
    .X(_09141_));
 sky130_fd_sc_hd__clkbuf_1 _14434_ (.A(_09141_),
    .X(_00345_));
 sky130_fd_sc_hd__buf_8 _14435_ (.A(net100),
    .X(_09142_));
 sky130_fd_sc_hd__clkbuf_8 _14436_ (.A(_09142_),
    .X(_09143_));
 sky130_fd_sc_hd__mux2_1 _14437_ (.A0(_09143_),
    .A1(net1679),
    .S(_09134_),
    .X(_09144_));
 sky130_fd_sc_hd__clkbuf_1 _14438_ (.A(_09144_),
    .X(_00346_));
 sky130_fd_sc_hd__buf_8 _14439_ (.A(net101),
    .X(_09145_));
 sky130_fd_sc_hd__buf_4 _14440_ (.A(_09145_),
    .X(_09146_));
 sky130_fd_sc_hd__mux2_1 _14441_ (.A0(_09146_),
    .A1(net996),
    .S(_09134_),
    .X(_09147_));
 sky130_fd_sc_hd__clkbuf_1 _14442_ (.A(_09147_),
    .X(_00347_));
 sky130_fd_sc_hd__buf_8 _14443_ (.A(net102),
    .X(_09148_));
 sky130_fd_sc_hd__buf_4 _14444_ (.A(_09148_),
    .X(_09149_));
 sky130_fd_sc_hd__mux2_1 _14445_ (.A0(_09149_),
    .A1(net841),
    .S(_09134_),
    .X(_09150_));
 sky130_fd_sc_hd__clkbuf_1 _14446_ (.A(_09150_),
    .X(_00348_));
 sky130_fd_sc_hd__buf_8 _14447_ (.A(net103),
    .X(_09151_));
 sky130_fd_sc_hd__buf_2 _14448_ (.A(_09151_),
    .X(_09152_));
 sky130_fd_sc_hd__mux2_1 _14449_ (.A0(_09152_),
    .A1(\cur_mb_mem[24][6] ),
    .S(_09134_),
    .X(_09153_));
 sky130_fd_sc_hd__clkbuf_1 _14450_ (.A(_09153_),
    .X(_00349_));
 sky130_fd_sc_hd__buf_8 _14451_ (.A(net104),
    .X(_09154_));
 sky130_fd_sc_hd__buf_4 _14452_ (.A(_09154_),
    .X(_09155_));
 sky130_fd_sc_hd__mux2_1 _14453_ (.A0(_09155_),
    .A1(\cur_mb_mem[24][7] ),
    .S(_09134_),
    .X(_09156_));
 sky130_fd_sc_hd__clkbuf_1 _14454_ (.A(_09156_),
    .X(_00350_));
 sky130_fd_sc_hd__nand2_8 _14455_ (.A(_06489_),
    .B(_09085_),
    .Y(_09157_));
 sky130_fd_sc_hd__mux2_1 _14456_ (.A0(_09133_),
    .A1(\cur_mb_mem[25][0] ),
    .S(_09157_),
    .X(_09158_));
 sky130_fd_sc_hd__clkbuf_1 _14457_ (.A(_09158_),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _14458_ (.A0(_09137_),
    .A1(net1828),
    .S(_09157_),
    .X(_09159_));
 sky130_fd_sc_hd__clkbuf_1 _14459_ (.A(_09159_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _14460_ (.A0(_09140_),
    .A1(net1936),
    .S(_09157_),
    .X(_09160_));
 sky130_fd_sc_hd__clkbuf_1 _14461_ (.A(_09160_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _14462_ (.A0(_09143_),
    .A1(\cur_mb_mem[25][3] ),
    .S(_09157_),
    .X(_09161_));
 sky130_fd_sc_hd__clkbuf_1 _14463_ (.A(_09161_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _14464_ (.A0(_09146_),
    .A1(net1531),
    .S(_09157_),
    .X(_09162_));
 sky130_fd_sc_hd__clkbuf_1 _14465_ (.A(_09162_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _14466_ (.A0(_09149_),
    .A1(net1377),
    .S(_09157_),
    .X(_09163_));
 sky130_fd_sc_hd__clkbuf_1 _14467_ (.A(_09163_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _14468_ (.A0(_09152_),
    .A1(\cur_mb_mem[25][6] ),
    .S(_09157_),
    .X(_09164_));
 sky130_fd_sc_hd__clkbuf_1 _14469_ (.A(_09164_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _14470_ (.A0(_09155_),
    .A1(\cur_mb_mem[25][7] ),
    .S(_09157_),
    .X(_09165_));
 sky130_fd_sc_hd__clkbuf_1 _14471_ (.A(_09165_),
    .X(_00358_));
 sky130_fd_sc_hd__nand2_8 _14472_ (.A(_06449_),
    .B(_09085_),
    .Y(_09166_));
 sky130_fd_sc_hd__mux2_1 _14473_ (.A0(_09133_),
    .A1(net1505),
    .S(_09166_),
    .X(_09167_));
 sky130_fd_sc_hd__clkbuf_1 _14474_ (.A(_09167_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _14475_ (.A0(_09137_),
    .A1(\cur_mb_mem[26][1] ),
    .S(_09166_),
    .X(_09168_));
 sky130_fd_sc_hd__clkbuf_1 _14476_ (.A(_09168_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _14477_ (.A0(_09140_),
    .A1(net1873),
    .S(_09166_),
    .X(_09169_));
 sky130_fd_sc_hd__clkbuf_1 _14478_ (.A(_09169_),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _14479_ (.A0(_09143_),
    .A1(\cur_mb_mem[26][3] ),
    .S(_09166_),
    .X(_09170_));
 sky130_fd_sc_hd__clkbuf_1 _14480_ (.A(_09170_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _14481_ (.A0(_09146_),
    .A1(net1752),
    .S(_09166_),
    .X(_09171_));
 sky130_fd_sc_hd__clkbuf_1 _14482_ (.A(_09171_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _14483_ (.A0(_09149_),
    .A1(net1768),
    .S(_09166_),
    .X(_09172_));
 sky130_fd_sc_hd__clkbuf_1 _14484_ (.A(_09172_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _14485_ (.A0(_09152_),
    .A1(net1647),
    .S(_09166_),
    .X(_09173_));
 sky130_fd_sc_hd__clkbuf_1 _14486_ (.A(_09173_),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _14487_ (.A0(_09155_),
    .A1(\cur_mb_mem[26][7] ),
    .S(_09166_),
    .X(_09174_));
 sky130_fd_sc_hd__clkbuf_1 _14488_ (.A(_09174_),
    .X(_00366_));
 sky130_fd_sc_hd__nand2_8 _14489_ (.A(_06476_),
    .B(_09085_),
    .Y(_09175_));
 sky130_fd_sc_hd__mux2_1 _14490_ (.A0(_09133_),
    .A1(net1788),
    .S(_09175_),
    .X(_09176_));
 sky130_fd_sc_hd__clkbuf_1 _14491_ (.A(_09176_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _14492_ (.A0(_09137_),
    .A1(\cur_mb_mem[27][1] ),
    .S(_09175_),
    .X(_09177_));
 sky130_fd_sc_hd__clkbuf_1 _14493_ (.A(_09177_),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _14494_ (.A0(_09140_),
    .A1(\cur_mb_mem[27][2] ),
    .S(_09175_),
    .X(_09178_));
 sky130_fd_sc_hd__clkbuf_1 _14495_ (.A(_09178_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _14496_ (.A0(_09143_),
    .A1(net612),
    .S(_09175_),
    .X(_09179_));
 sky130_fd_sc_hd__clkbuf_1 _14497_ (.A(_09179_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _14498_ (.A0(_09146_),
    .A1(net1568),
    .S(_09175_),
    .X(_09180_));
 sky130_fd_sc_hd__clkbuf_1 _14499_ (.A(_09180_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _14500_ (.A0(_09149_),
    .A1(net1670),
    .S(_09175_),
    .X(_09181_));
 sky130_fd_sc_hd__clkbuf_1 _14501_ (.A(_09181_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _14502_ (.A0(_09152_),
    .A1(net1906),
    .S(_09175_),
    .X(_09182_));
 sky130_fd_sc_hd__clkbuf_1 _14503_ (.A(_09182_),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _14504_ (.A0(_09155_),
    .A1(\cur_mb_mem[27][7] ),
    .S(_09175_),
    .X(_09183_));
 sky130_fd_sc_hd__clkbuf_1 _14505_ (.A(_09183_),
    .X(_00374_));
 sky130_fd_sc_hd__nand2_8 _14506_ (.A(_06017_),
    .B(_09085_),
    .Y(_09184_));
 sky130_fd_sc_hd__mux2_1 _14507_ (.A0(_09133_),
    .A1(net1698),
    .S(_09184_),
    .X(_09185_));
 sky130_fd_sc_hd__clkbuf_1 _14508_ (.A(_09185_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _14509_ (.A0(_09137_),
    .A1(\cur_mb_mem[28][1] ),
    .S(_09184_),
    .X(_09186_));
 sky130_fd_sc_hd__clkbuf_1 _14510_ (.A(_09186_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _14511_ (.A0(_09140_),
    .A1(net1614),
    .S(_09184_),
    .X(_09187_));
 sky130_fd_sc_hd__clkbuf_1 _14512_ (.A(_09187_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _14513_ (.A0(_09143_),
    .A1(\cur_mb_mem[28][3] ),
    .S(_09184_),
    .X(_09188_));
 sky130_fd_sc_hd__clkbuf_1 _14514_ (.A(_09188_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _14515_ (.A0(_09146_),
    .A1(net1732),
    .S(_09184_),
    .X(_09189_));
 sky130_fd_sc_hd__clkbuf_1 _14516_ (.A(_09189_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _14517_ (.A0(_09149_),
    .A1(net951),
    .S(_09184_),
    .X(_09190_));
 sky130_fd_sc_hd__clkbuf_1 _14518_ (.A(_09190_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _14519_ (.A0(_09152_),
    .A1(net1457),
    .S(_09184_),
    .X(_09191_));
 sky130_fd_sc_hd__clkbuf_1 _14520_ (.A(_09191_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _14521_ (.A0(_09155_),
    .A1(\cur_mb_mem[28][7] ),
    .S(_09184_),
    .X(_09192_));
 sky130_fd_sc_hd__clkbuf_1 _14522_ (.A(_09192_),
    .X(_00382_));
 sky130_fd_sc_hd__nand2_8 _14523_ (.A(_06404_),
    .B(_09085_),
    .Y(_09193_));
 sky130_fd_sc_hd__mux2_1 _14524_ (.A0(_09133_),
    .A1(net1657),
    .S(_09193_),
    .X(_09194_));
 sky130_fd_sc_hd__clkbuf_1 _14525_ (.A(_09194_),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _14526_ (.A0(_09137_),
    .A1(\cur_mb_mem[29][1] ),
    .S(_09193_),
    .X(_09195_));
 sky130_fd_sc_hd__clkbuf_1 _14527_ (.A(_09195_),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _14528_ (.A0(_09140_),
    .A1(net1803),
    .S(_09193_),
    .X(_09196_));
 sky130_fd_sc_hd__clkbuf_1 _14529_ (.A(_09196_),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _14530_ (.A0(_09143_),
    .A1(net1926),
    .S(_09193_),
    .X(_09197_));
 sky130_fd_sc_hd__clkbuf_1 _14531_ (.A(_09197_),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _14532_ (.A0(_09146_),
    .A1(net1515),
    .S(_09193_),
    .X(_09198_));
 sky130_fd_sc_hd__clkbuf_1 _14533_ (.A(_09198_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _14534_ (.A0(_09149_),
    .A1(net1555),
    .S(_09193_),
    .X(_09199_));
 sky130_fd_sc_hd__clkbuf_1 _14535_ (.A(_09199_),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _14536_ (.A0(_09152_),
    .A1(\cur_mb_mem[29][6] ),
    .S(_09193_),
    .X(_09200_));
 sky130_fd_sc_hd__clkbuf_1 _14537_ (.A(_09200_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _14538_ (.A0(_09155_),
    .A1(\cur_mb_mem[29][7] ),
    .S(_09193_),
    .X(_09201_));
 sky130_fd_sc_hd__clkbuf_1 _14539_ (.A(_09201_),
    .X(_00390_));
 sky130_fd_sc_hd__nand2_8 _14540_ (.A(_06002_),
    .B(_09085_),
    .Y(_09202_));
 sky130_fd_sc_hd__mux2_1 _14541_ (.A0(_09133_),
    .A1(net1414),
    .S(_09202_),
    .X(_09203_));
 sky130_fd_sc_hd__clkbuf_1 _14542_ (.A(_09203_),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _14543_ (.A0(_09137_),
    .A1(net973),
    .S(_09202_),
    .X(_09204_));
 sky130_fd_sc_hd__clkbuf_1 _14544_ (.A(_09204_),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _14545_ (.A0(_09140_),
    .A1(net1760),
    .S(_09202_),
    .X(_09205_));
 sky130_fd_sc_hd__clkbuf_1 _14546_ (.A(_09205_),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _14547_ (.A0(_09143_),
    .A1(net1758),
    .S(_09202_),
    .X(_09206_));
 sky130_fd_sc_hd__clkbuf_1 _14548_ (.A(_09206_),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _14549_ (.A0(_09146_),
    .A1(net1573),
    .S(_09202_),
    .X(_09207_));
 sky130_fd_sc_hd__clkbuf_1 _14550_ (.A(_09207_),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _14551_ (.A0(_09149_),
    .A1(net1635),
    .S(_09202_),
    .X(_09208_));
 sky130_fd_sc_hd__clkbuf_1 _14552_ (.A(_09208_),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _14553_ (.A0(_09152_),
    .A1(net1946),
    .S(_09202_),
    .X(_09209_));
 sky130_fd_sc_hd__clkbuf_1 _14554_ (.A(_09209_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _14555_ (.A0(_09155_),
    .A1(\cur_mb_mem[30][7] ),
    .S(_09202_),
    .X(_09210_));
 sky130_fd_sc_hd__clkbuf_1 _14556_ (.A(_09210_),
    .X(_00398_));
 sky130_fd_sc_hd__buf_12 _14557_ (.A(_08901_),
    .X(_09211_));
 sky130_fd_sc_hd__nand2_8 _14558_ (.A(_06178_),
    .B(_09211_),
    .Y(_09212_));
 sky130_fd_sc_hd__mux2_1 _14559_ (.A0(_09133_),
    .A1(net1456),
    .S(_09212_),
    .X(_09213_));
 sky130_fd_sc_hd__clkbuf_1 _14560_ (.A(_09213_),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _14561_ (.A0(_09137_),
    .A1(\cur_mb_mem[31][1] ),
    .S(_09212_),
    .X(_09214_));
 sky130_fd_sc_hd__clkbuf_1 _14562_ (.A(_09214_),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _14563_ (.A0(_09140_),
    .A1(net1987),
    .S(_09212_),
    .X(_09215_));
 sky130_fd_sc_hd__clkbuf_1 _14564_ (.A(_09215_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _14565_ (.A0(_09143_),
    .A1(net1799),
    .S(_09212_),
    .X(_09216_));
 sky130_fd_sc_hd__clkbuf_1 _14566_ (.A(_09216_),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _14567_ (.A0(_09146_),
    .A1(net1903),
    .S(_09212_),
    .X(_09217_));
 sky130_fd_sc_hd__clkbuf_1 _14568_ (.A(_09217_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _14569_ (.A0(_09149_),
    .A1(net1834),
    .S(_09212_),
    .X(_09218_));
 sky130_fd_sc_hd__clkbuf_1 _14570_ (.A(_09218_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _14571_ (.A0(_09152_),
    .A1(\cur_mb_mem[31][6] ),
    .S(_09212_),
    .X(_09219_));
 sky130_fd_sc_hd__clkbuf_1 _14572_ (.A(_09219_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _14573_ (.A0(_09155_),
    .A1(\cur_mb_mem[31][7] ),
    .S(_09212_),
    .X(_09220_));
 sky130_fd_sc_hd__clkbuf_1 _14574_ (.A(_09220_),
    .X(_00406_));
 sky130_fd_sc_hd__nand2_8 _14575_ (.A(_06044_),
    .B(_08883_),
    .Y(_09221_));
 sky130_fd_sc_hd__mux2_1 _14576_ (.A0(_09133_),
    .A1(net1539),
    .S(_09221_),
    .X(_09222_));
 sky130_fd_sc_hd__clkbuf_1 _14577_ (.A(_09222_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _14578_ (.A0(_09137_),
    .A1(\cur_mb_mem[32][1] ),
    .S(_09221_),
    .X(_09223_));
 sky130_fd_sc_hd__clkbuf_1 _14579_ (.A(_09223_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _14580_ (.A0(_09140_),
    .A1(\cur_mb_mem[32][2] ),
    .S(_09221_),
    .X(_09224_));
 sky130_fd_sc_hd__clkbuf_1 _14581_ (.A(_09224_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _14582_ (.A0(_09143_),
    .A1(net1992),
    .S(_09221_),
    .X(_09225_));
 sky130_fd_sc_hd__clkbuf_1 _14583_ (.A(_09225_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _14584_ (.A0(_09146_),
    .A1(net1928),
    .S(_09221_),
    .X(_09226_));
 sky130_fd_sc_hd__clkbuf_1 _14585_ (.A(_09226_),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _14586_ (.A0(_09149_),
    .A1(net1895),
    .S(_09221_),
    .X(_09227_));
 sky130_fd_sc_hd__clkbuf_1 _14587_ (.A(_09227_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _14588_ (.A0(_09152_),
    .A1(\cur_mb_mem[32][6] ),
    .S(_09221_),
    .X(_09228_));
 sky130_fd_sc_hd__clkbuf_1 _14589_ (.A(_09228_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _14590_ (.A0(_09155_),
    .A1(\cur_mb_mem[32][7] ),
    .S(_09221_),
    .X(_09229_));
 sky130_fd_sc_hd__clkbuf_1 _14591_ (.A(_09229_),
    .X(_00414_));
 sky130_fd_sc_hd__nand2_8 _14592_ (.A(_06291_),
    .B(_09211_),
    .Y(_09230_));
 sky130_fd_sc_hd__mux2_1 _14593_ (.A0(_09133_),
    .A1(\cur_mb_mem[33][0] ),
    .S(_09230_),
    .X(_09231_));
 sky130_fd_sc_hd__clkbuf_1 _14594_ (.A(_09231_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _14595_ (.A0(_09137_),
    .A1(net1704),
    .S(_09230_),
    .X(_09232_));
 sky130_fd_sc_hd__clkbuf_1 _14596_ (.A(_09232_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _14597_ (.A0(_09140_),
    .A1(\cur_mb_mem[33][2] ),
    .S(_09230_),
    .X(_09233_));
 sky130_fd_sc_hd__clkbuf_1 _14598_ (.A(_09233_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _14599_ (.A0(_09143_),
    .A1(net511),
    .S(_09230_),
    .X(_09234_));
 sky130_fd_sc_hd__clkbuf_1 _14600_ (.A(_09234_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _14601_ (.A0(_09146_),
    .A1(\cur_mb_mem[33][4] ),
    .S(_09230_),
    .X(_09235_));
 sky130_fd_sc_hd__clkbuf_1 _14602_ (.A(_09235_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _14603_ (.A0(_09149_),
    .A1(\cur_mb_mem[33][5] ),
    .S(_09230_),
    .X(_09236_));
 sky130_fd_sc_hd__clkbuf_1 _14604_ (.A(_09236_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _14605_ (.A0(_09152_),
    .A1(net1925),
    .S(_09230_),
    .X(_09237_));
 sky130_fd_sc_hd__clkbuf_1 _14606_ (.A(_09237_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _14607_ (.A0(_09155_),
    .A1(net1153),
    .S(_09230_),
    .X(_09238_));
 sky130_fd_sc_hd__clkbuf_1 _14608_ (.A(_09238_),
    .X(_00422_));
 sky130_fd_sc_hd__buf_8 _14609_ (.A(_09132_),
    .X(_09239_));
 sky130_fd_sc_hd__nand2_8 _14610_ (.A(_06393_),
    .B(_09211_),
    .Y(_09240_));
 sky130_fd_sc_hd__mux2_1 _14611_ (.A0(_09239_),
    .A1(net738),
    .S(_09240_),
    .X(_09241_));
 sky130_fd_sc_hd__clkbuf_1 _14612_ (.A(_09241_),
    .X(_00423_));
 sky130_fd_sc_hd__buf_8 _14613_ (.A(_09136_),
    .X(_09242_));
 sky130_fd_sc_hd__mux2_1 _14614_ (.A0(_09242_),
    .A1(net1331),
    .S(_09240_),
    .X(_09243_));
 sky130_fd_sc_hd__clkbuf_1 _14615_ (.A(_09243_),
    .X(_00424_));
 sky130_fd_sc_hd__buf_8 _14616_ (.A(_09139_),
    .X(_09244_));
 sky130_fd_sc_hd__mux2_1 _14617_ (.A0(_09244_),
    .A1(net1044),
    .S(_09240_),
    .X(_09245_));
 sky130_fd_sc_hd__clkbuf_1 _14618_ (.A(_09245_),
    .X(_00425_));
 sky130_fd_sc_hd__buf_8 _14619_ (.A(_09142_),
    .X(_09246_));
 sky130_fd_sc_hd__mux2_1 _14620_ (.A0(_09246_),
    .A1(net626),
    .S(_09240_),
    .X(_09247_));
 sky130_fd_sc_hd__clkbuf_1 _14621_ (.A(_09247_),
    .X(_00426_));
 sky130_fd_sc_hd__clkbuf_16 _14622_ (.A(_09145_),
    .X(_09248_));
 sky130_fd_sc_hd__mux2_1 _14623_ (.A0(_09248_),
    .A1(net1172),
    .S(_09240_),
    .X(_09249_));
 sky130_fd_sc_hd__clkbuf_1 _14624_ (.A(_09249_),
    .X(_00427_));
 sky130_fd_sc_hd__clkbuf_16 _14625_ (.A(_09148_),
    .X(_09250_));
 sky130_fd_sc_hd__mux2_1 _14626_ (.A0(_09250_),
    .A1(net1283),
    .S(_09240_),
    .X(_09251_));
 sky130_fd_sc_hd__clkbuf_1 _14627_ (.A(_09251_),
    .X(_00428_));
 sky130_fd_sc_hd__buf_6 _14628_ (.A(_09151_),
    .X(_09252_));
 sky130_fd_sc_hd__mux2_1 _14629_ (.A0(_09252_),
    .A1(net1193),
    .S(_09240_),
    .X(_09253_));
 sky130_fd_sc_hd__clkbuf_1 _14630_ (.A(_09253_),
    .X(_00429_));
 sky130_fd_sc_hd__buf_6 _14631_ (.A(_09154_),
    .X(_09254_));
 sky130_fd_sc_hd__mux2_1 _14632_ (.A0(_09254_),
    .A1(net1224),
    .S(_09240_),
    .X(_09255_));
 sky130_fd_sc_hd__clkbuf_1 _14633_ (.A(_09255_),
    .X(_00430_));
 sky130_fd_sc_hd__nand2_8 _14634_ (.A(_06088_),
    .B(_09211_),
    .Y(_09256_));
 sky130_fd_sc_hd__mux2_1 _14635_ (.A0(_09239_),
    .A1(net978),
    .S(_09256_),
    .X(_09257_));
 sky130_fd_sc_hd__clkbuf_1 _14636_ (.A(_09257_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _14637_ (.A0(_09242_),
    .A1(\cur_mb_mem[35][1] ),
    .S(_09256_),
    .X(_09258_));
 sky130_fd_sc_hd__clkbuf_1 _14638_ (.A(_09258_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _14639_ (.A0(_09244_),
    .A1(net1811),
    .S(_09256_),
    .X(_09259_));
 sky130_fd_sc_hd__clkbuf_1 _14640_ (.A(_09259_),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _14641_ (.A0(_09246_),
    .A1(net1010),
    .S(_09256_),
    .X(_09260_));
 sky130_fd_sc_hd__clkbuf_1 _14642_ (.A(_09260_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _14643_ (.A0(_09248_),
    .A1(net718),
    .S(_09256_),
    .X(_09261_));
 sky130_fd_sc_hd__clkbuf_1 _14644_ (.A(_09261_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _14645_ (.A0(_09250_),
    .A1(net799),
    .S(_09256_),
    .X(_09262_));
 sky130_fd_sc_hd__clkbuf_1 _14646_ (.A(_09262_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _14647_ (.A0(_09252_),
    .A1(net1547),
    .S(_09256_),
    .X(_09263_));
 sky130_fd_sc_hd__clkbuf_1 _14648_ (.A(_09263_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _14649_ (.A0(_09254_),
    .A1(net1209),
    .S(_09256_),
    .X(_09264_));
 sky130_fd_sc_hd__clkbuf_1 _14650_ (.A(_09264_),
    .X(_00438_));
 sky130_fd_sc_hd__nand2_8 _14651_ (.A(_06360_),
    .B(_09211_),
    .Y(_09265_));
 sky130_fd_sc_hd__mux2_1 _14652_ (.A0(_09239_),
    .A1(net1318),
    .S(_09265_),
    .X(_09266_));
 sky130_fd_sc_hd__clkbuf_1 _14653_ (.A(_09266_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _14654_ (.A0(_09242_),
    .A1(net1749),
    .S(_09265_),
    .X(_09267_));
 sky130_fd_sc_hd__clkbuf_1 _14655_ (.A(_09267_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _14656_ (.A0(_09244_),
    .A1(net1175),
    .S(_09265_),
    .X(_09268_));
 sky130_fd_sc_hd__clkbuf_1 _14657_ (.A(_09268_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _14658_ (.A0(_09246_),
    .A1(net1188),
    .S(_09265_),
    .X(_09269_));
 sky130_fd_sc_hd__clkbuf_1 _14659_ (.A(_09269_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _14660_ (.A0(_09248_),
    .A1(net898),
    .S(_09265_),
    .X(_09270_));
 sky130_fd_sc_hd__clkbuf_1 _14661_ (.A(_09270_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _14662_ (.A0(_09250_),
    .A1(net701),
    .S(_09265_),
    .X(_09271_));
 sky130_fd_sc_hd__clkbuf_1 _14663_ (.A(_09271_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _14664_ (.A0(_09252_),
    .A1(net1466),
    .S(_09265_),
    .X(_09272_));
 sky130_fd_sc_hd__clkbuf_1 _14665_ (.A(_09272_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _14666_ (.A0(_09254_),
    .A1(net1144),
    .S(_09265_),
    .X(_09273_));
 sky130_fd_sc_hd__clkbuf_1 _14667_ (.A(_09273_),
    .X(_00446_));
 sky130_fd_sc_hd__nand2_4 _14668_ (.A(_06344_),
    .B(_09211_),
    .Y(_09274_));
 sky130_fd_sc_hd__mux2_1 _14669_ (.A0(_09239_),
    .A1(net1092),
    .S(_09274_),
    .X(_09275_));
 sky130_fd_sc_hd__clkbuf_1 _14670_ (.A(_09275_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _14671_ (.A0(_09242_),
    .A1(net1462),
    .S(_09274_),
    .X(_09276_));
 sky130_fd_sc_hd__clkbuf_1 _14672_ (.A(_09276_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _14673_ (.A0(_09244_),
    .A1(net1783),
    .S(_09274_),
    .X(_09277_));
 sky130_fd_sc_hd__clkbuf_1 _14674_ (.A(_09277_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _14675_ (.A0(_09246_),
    .A1(net1418),
    .S(_09274_),
    .X(_09278_));
 sky130_fd_sc_hd__clkbuf_1 _14676_ (.A(_09278_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _14677_ (.A0(_09248_),
    .A1(net601),
    .S(_09274_),
    .X(_09279_));
 sky130_fd_sc_hd__clkbuf_1 _14678_ (.A(_09279_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _14679_ (.A0(_09250_),
    .A1(net882),
    .S(_09274_),
    .X(_09280_));
 sky130_fd_sc_hd__clkbuf_1 _14680_ (.A(_09280_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _14681_ (.A0(_09252_),
    .A1(net1500),
    .S(_09274_),
    .X(_09281_));
 sky130_fd_sc_hd__clkbuf_1 _14682_ (.A(_09281_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _14683_ (.A0(_09254_),
    .A1(net1221),
    .S(_09274_),
    .X(_09282_));
 sky130_fd_sc_hd__clkbuf_1 _14684_ (.A(_09282_),
    .X(_00454_));
 sky130_fd_sc_hd__nand2_8 _14685_ (.A(_06396_),
    .B(_09211_),
    .Y(_09283_));
 sky130_fd_sc_hd__mux2_1 _14686_ (.A0(_09239_),
    .A1(net1536),
    .S(_09283_),
    .X(_09284_));
 sky130_fd_sc_hd__clkbuf_1 _14687_ (.A(_09284_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _14688_ (.A0(_09242_),
    .A1(net1233),
    .S(_09283_),
    .X(_09285_));
 sky130_fd_sc_hd__clkbuf_1 _14689_ (.A(_09285_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _14690_ (.A0(_09244_),
    .A1(net1559),
    .S(_09283_),
    .X(_09286_));
 sky130_fd_sc_hd__clkbuf_1 _14691_ (.A(_09286_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _14692_ (.A0(_09246_),
    .A1(net1488),
    .S(_09283_),
    .X(_09287_));
 sky130_fd_sc_hd__clkbuf_1 _14693_ (.A(_09287_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _14694_ (.A0(_09248_),
    .A1(net1286),
    .S(_09283_),
    .X(_09288_));
 sky130_fd_sc_hd__clkbuf_1 _14695_ (.A(_09288_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _14696_ (.A0(_09250_),
    .A1(net1397),
    .S(_09283_),
    .X(_09289_));
 sky130_fd_sc_hd__clkbuf_1 _14697_ (.A(_09289_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _14698_ (.A0(_09252_),
    .A1(\cur_mb_mem[38][6] ),
    .S(_09283_),
    .X(_09290_));
 sky130_fd_sc_hd__clkbuf_1 _14699_ (.A(_09290_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _14700_ (.A0(_09254_),
    .A1(net1994),
    .S(_09283_),
    .X(_09291_));
 sky130_fd_sc_hd__clkbuf_1 _14701_ (.A(_09291_),
    .X(_00462_));
 sky130_fd_sc_hd__nand2_4 _14702_ (.A(_06373_),
    .B(_09211_),
    .Y(_09292_));
 sky130_fd_sc_hd__mux2_1 _14703_ (.A0(_09239_),
    .A1(net1360),
    .S(_09292_),
    .X(_09293_));
 sky130_fd_sc_hd__clkbuf_1 _14704_ (.A(_09293_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _14705_ (.A0(_09242_),
    .A1(net546),
    .S(_09292_),
    .X(_09294_));
 sky130_fd_sc_hd__clkbuf_1 _14706_ (.A(_09294_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _14707_ (.A0(_09244_),
    .A1(net1644),
    .S(_09292_),
    .X(_09295_));
 sky130_fd_sc_hd__clkbuf_1 _14708_ (.A(_09295_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _14709_ (.A0(_09246_),
    .A1(net1315),
    .S(_09292_),
    .X(_09296_));
 sky130_fd_sc_hd__clkbuf_1 _14710_ (.A(_09296_),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _14711_ (.A0(_09248_),
    .A1(net805),
    .S(_09292_),
    .X(_09297_));
 sky130_fd_sc_hd__clkbuf_1 _14712_ (.A(_09297_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _14713_ (.A0(_09250_),
    .A1(net1099),
    .S(_09292_),
    .X(_09298_));
 sky130_fd_sc_hd__clkbuf_1 _14714_ (.A(_09298_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _14715_ (.A0(_09252_),
    .A1(net1571),
    .S(_09292_),
    .X(_09299_));
 sky130_fd_sc_hd__clkbuf_1 _14716_ (.A(_09299_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _14717_ (.A0(_09254_),
    .A1(net1910),
    .S(_09292_),
    .X(_09300_));
 sky130_fd_sc_hd__clkbuf_1 _14718_ (.A(_09300_),
    .X(_00470_));
 sky130_fd_sc_hd__nand2_8 _14719_ (.A(_06485_),
    .B(_09211_),
    .Y(_09301_));
 sky130_fd_sc_hd__mux2_1 _14720_ (.A0(_09239_),
    .A1(net663),
    .S(_09301_),
    .X(_09302_));
 sky130_fd_sc_hd__clkbuf_1 _14721_ (.A(_09302_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _14722_ (.A0(_09242_),
    .A1(net1191),
    .S(_09301_),
    .X(_09303_));
 sky130_fd_sc_hd__clkbuf_1 _14723_ (.A(_09303_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _14724_ (.A0(_09244_),
    .A1(net992),
    .S(_09301_),
    .X(_09304_));
 sky130_fd_sc_hd__clkbuf_1 _14725_ (.A(_09304_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _14726_ (.A0(_09246_),
    .A1(net806),
    .S(_09301_),
    .X(_09305_));
 sky130_fd_sc_hd__clkbuf_1 _14727_ (.A(_09305_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _14728_ (.A0(_09248_),
    .A1(net1415),
    .S(_09301_),
    .X(_09306_));
 sky130_fd_sc_hd__clkbuf_1 _14729_ (.A(_09306_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _14730_ (.A0(_09250_),
    .A1(net1592),
    .S(_09301_),
    .X(_09307_));
 sky130_fd_sc_hd__clkbuf_1 _14731_ (.A(_09307_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _14732_ (.A0(_09252_),
    .A1(net1398),
    .S(_09301_),
    .X(_09308_));
 sky130_fd_sc_hd__clkbuf_1 _14733_ (.A(_09308_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _14734_ (.A0(_09254_),
    .A1(net1575),
    .S(_09301_),
    .X(_09309_));
 sky130_fd_sc_hd__clkbuf_1 _14735_ (.A(_09309_),
    .X(_00478_));
 sky130_fd_sc_hd__nand2_8 _14736_ (.A(_06031_),
    .B(_09211_),
    .Y(_09310_));
 sky130_fd_sc_hd__mux2_1 _14737_ (.A0(_09239_),
    .A1(net870),
    .S(_09310_),
    .X(_09311_));
 sky130_fd_sc_hd__clkbuf_1 _14738_ (.A(_09311_),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _14739_ (.A0(_09242_),
    .A1(net1616),
    .S(_09310_),
    .X(_09312_));
 sky130_fd_sc_hd__clkbuf_1 _14740_ (.A(_09312_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _14741_ (.A0(_09244_),
    .A1(net775),
    .S(_09310_),
    .X(_09313_));
 sky130_fd_sc_hd__clkbuf_1 _14742_ (.A(_09313_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _14743_ (.A0(_09246_),
    .A1(net1490),
    .S(_09310_),
    .X(_09314_));
 sky130_fd_sc_hd__clkbuf_1 _14744_ (.A(_09314_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _14745_ (.A0(_09248_),
    .A1(net1438),
    .S(_09310_),
    .X(_09315_));
 sky130_fd_sc_hd__clkbuf_1 _14746_ (.A(_09315_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _14747_ (.A0(_09250_),
    .A1(net1168),
    .S(_09310_),
    .X(_09316_));
 sky130_fd_sc_hd__clkbuf_1 _14748_ (.A(_09316_),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _14749_ (.A0(_09252_),
    .A1(\cur_mb_mem[41][6] ),
    .S(_09310_),
    .X(_09317_));
 sky130_fd_sc_hd__clkbuf_1 _14750_ (.A(_09317_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _14751_ (.A0(_09254_),
    .A1(net1136),
    .S(_09310_),
    .X(_09318_));
 sky130_fd_sc_hd__clkbuf_1 _14752_ (.A(_09318_),
    .X(_00486_));
 sky130_fd_sc_hd__buf_12 _14753_ (.A(_08958_),
    .X(_09319_));
 sky130_fd_sc_hd__nand2_8 _14754_ (.A(_06441_),
    .B(_09319_),
    .Y(_09320_));
 sky130_fd_sc_hd__mux2_1 _14755_ (.A0(_09239_),
    .A1(net1535),
    .S(_09320_),
    .X(_09321_));
 sky130_fd_sc_hd__clkbuf_1 _14756_ (.A(_09321_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _14757_ (.A0(_09242_),
    .A1(\cur_mb_mem[42][1] ),
    .S(_09320_),
    .X(_09322_));
 sky130_fd_sc_hd__clkbuf_1 _14758_ (.A(_09322_),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _14759_ (.A0(_09244_),
    .A1(net1150),
    .S(_09320_),
    .X(_09323_));
 sky130_fd_sc_hd__clkbuf_1 _14760_ (.A(_09323_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _14761_ (.A0(_09246_),
    .A1(net1229),
    .S(_09320_),
    .X(_09324_));
 sky130_fd_sc_hd__clkbuf_1 _14762_ (.A(_09324_),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _14763_ (.A0(_09248_),
    .A1(net1423),
    .S(_09320_),
    .X(_09325_));
 sky130_fd_sc_hd__clkbuf_1 _14764_ (.A(_09325_),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _14765_ (.A0(_09250_),
    .A1(net1164),
    .S(_09320_),
    .X(_09326_));
 sky130_fd_sc_hd__clkbuf_1 _14766_ (.A(_09326_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _14767_ (.A0(_09252_),
    .A1(net1309),
    .S(_09320_),
    .X(_09327_));
 sky130_fd_sc_hd__clkbuf_1 _14768_ (.A(_09327_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _14769_ (.A0(_09254_),
    .A1(net1684),
    .S(_09320_),
    .X(_09328_));
 sky130_fd_sc_hd__clkbuf_1 _14770_ (.A(_09328_),
    .X(_00494_));
 sky130_fd_sc_hd__nand2_8 _14771_ (.A(_06006_),
    .B(_09319_),
    .Y(_09329_));
 sky130_fd_sc_hd__mux2_1 _14772_ (.A0(_09239_),
    .A1(net576),
    .S(_09329_),
    .X(_09330_));
 sky130_fd_sc_hd__clkbuf_1 _14773_ (.A(_09330_),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _14774_ (.A0(_09242_),
    .A1(net1371),
    .S(_09329_),
    .X(_09331_));
 sky130_fd_sc_hd__clkbuf_1 _14775_ (.A(_09331_),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _14776_ (.A0(_09244_),
    .A1(net704),
    .S(_09329_),
    .X(_09332_));
 sky130_fd_sc_hd__clkbuf_1 _14777_ (.A(_09332_),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _14778_ (.A0(_09246_),
    .A1(net715),
    .S(_09329_),
    .X(_09333_));
 sky130_fd_sc_hd__clkbuf_1 _14779_ (.A(_09333_),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _14780_ (.A0(_09248_),
    .A1(net1432),
    .S(_09329_),
    .X(_09334_));
 sky130_fd_sc_hd__clkbuf_1 _14781_ (.A(_09334_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _14782_ (.A0(_09250_),
    .A1(net1155),
    .S(_09329_),
    .X(_02191_));
 sky130_fd_sc_hd__clkbuf_1 _14783_ (.A(_02191_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _14784_ (.A0(_09252_),
    .A1(net1314),
    .S(_09329_),
    .X(_02192_));
 sky130_fd_sc_hd__clkbuf_1 _14785_ (.A(_02192_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _14786_ (.A0(_09254_),
    .A1(net1542),
    .S(_09329_),
    .X(_02193_));
 sky130_fd_sc_hd__clkbuf_1 _14787_ (.A(_02193_),
    .X(_00502_));
 sky130_fd_sc_hd__buf_12 _14788_ (.A(_09132_),
    .X(_02194_));
 sky130_fd_sc_hd__nand2_8 _14789_ (.A(_06399_),
    .B(_09319_),
    .Y(_02195_));
 sky130_fd_sc_hd__mux2_1 _14790_ (.A0(_02194_),
    .A1(net1232),
    .S(_02195_),
    .X(_02196_));
 sky130_fd_sc_hd__clkbuf_1 _14791_ (.A(_02196_),
    .X(_00503_));
 sky130_fd_sc_hd__buf_4 _14792_ (.A(_09136_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _14793_ (.A0(_02197_),
    .A1(net1247),
    .S(_02195_),
    .X(_02198_));
 sky130_fd_sc_hd__clkbuf_1 _14794_ (.A(_02198_),
    .X(_00504_));
 sky130_fd_sc_hd__clkbuf_16 _14795_ (.A(_09139_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_1 _14796_ (.A0(_02199_),
    .A1(net1558),
    .S(_02195_),
    .X(_02200_));
 sky130_fd_sc_hd__clkbuf_1 _14797_ (.A(_02200_),
    .X(_00505_));
 sky130_fd_sc_hd__clkbuf_16 _14798_ (.A(_09142_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _14799_ (.A0(_02201_),
    .A1(net1277),
    .S(_02195_),
    .X(_02202_));
 sky130_fd_sc_hd__clkbuf_1 _14800_ (.A(_02202_),
    .X(_00506_));
 sky130_fd_sc_hd__clkbuf_8 _14801_ (.A(_09145_),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_1 _14802_ (.A0(_02203_),
    .A1(net947),
    .S(_02195_),
    .X(_02204_));
 sky130_fd_sc_hd__clkbuf_1 _14803_ (.A(_02204_),
    .X(_00507_));
 sky130_fd_sc_hd__clkbuf_8 _14804_ (.A(_09148_),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_1 _14805_ (.A0(_02205_),
    .A1(net764),
    .S(_02195_),
    .X(_02206_));
 sky130_fd_sc_hd__clkbuf_1 _14806_ (.A(_02206_),
    .X(_00508_));
 sky130_fd_sc_hd__buf_6 _14807_ (.A(_09151_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _14808_ (.A0(_02207_),
    .A1(net1428),
    .S(_02195_),
    .X(_02208_));
 sky130_fd_sc_hd__clkbuf_1 _14809_ (.A(_02208_),
    .X(_00509_));
 sky130_fd_sc_hd__buf_8 _14810_ (.A(_09154_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _14811_ (.A0(_02209_),
    .A1(net1449),
    .S(_02195_),
    .X(_02210_));
 sky130_fd_sc_hd__clkbuf_1 _14812_ (.A(_02210_),
    .X(_00510_));
 sky130_fd_sc_hd__nand2_8 _14813_ (.A(_06491_),
    .B(_09319_),
    .Y(_02211_));
 sky130_fd_sc_hd__mux2_1 _14814_ (.A0(_02194_),
    .A1(net1460),
    .S(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__clkbuf_1 _14815_ (.A(_02212_),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _14816_ (.A0(_02197_),
    .A1(\cur_mb_mem[45][1] ),
    .S(_02211_),
    .X(_02213_));
 sky130_fd_sc_hd__clkbuf_1 _14817_ (.A(_02213_),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _14818_ (.A0(_02199_),
    .A1(net1433),
    .S(_02211_),
    .X(_02214_));
 sky130_fd_sc_hd__clkbuf_1 _14819_ (.A(_02214_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _14820_ (.A0(_02201_),
    .A1(net1608),
    .S(_02211_),
    .X(_02215_));
 sky130_fd_sc_hd__clkbuf_1 _14821_ (.A(_02215_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _14822_ (.A0(_02203_),
    .A1(net1735),
    .S(_02211_),
    .X(_02216_));
 sky130_fd_sc_hd__clkbuf_1 _14823_ (.A(_02216_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _14824_ (.A0(_02205_),
    .A1(net1791),
    .S(_02211_),
    .X(_02217_));
 sky130_fd_sc_hd__clkbuf_1 _14825_ (.A(_02217_),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _14826_ (.A0(_02207_),
    .A1(net1622),
    .S(_02211_),
    .X(_02218_));
 sky130_fd_sc_hd__clkbuf_1 _14827_ (.A(_02218_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _14828_ (.A0(_02209_),
    .A1(net1708),
    .S(_02211_),
    .X(_02219_));
 sky130_fd_sc_hd__clkbuf_1 _14829_ (.A(_02219_),
    .X(_00518_));
 sky130_fd_sc_hd__nand2_8 _14830_ (.A(_06107_),
    .B(_09319_),
    .Y(_02220_));
 sky130_fd_sc_hd__mux2_1 _14831_ (.A0(_02194_),
    .A1(net867),
    .S(_02220_),
    .X(_02221_));
 sky130_fd_sc_hd__clkbuf_1 _14832_ (.A(_02221_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _14833_ (.A0(_02197_),
    .A1(net1196),
    .S(_02220_),
    .X(_02222_));
 sky130_fd_sc_hd__clkbuf_1 _14834_ (.A(_02222_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _14835_ (.A0(_02199_),
    .A1(net1454),
    .S(_02220_),
    .X(_02223_));
 sky130_fd_sc_hd__clkbuf_1 _14836_ (.A(_02223_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _14837_ (.A0(_02201_),
    .A1(net1386),
    .S(_02220_),
    .X(_02224_));
 sky130_fd_sc_hd__clkbuf_1 _14838_ (.A(_02224_),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _14839_ (.A0(_02203_),
    .A1(net960),
    .S(_02220_),
    .X(_02225_));
 sky130_fd_sc_hd__clkbuf_1 _14840_ (.A(_02225_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _14841_ (.A0(_02205_),
    .A1(net1308),
    .S(_02220_),
    .X(_02226_));
 sky130_fd_sc_hd__clkbuf_1 _14842_ (.A(_02226_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _14843_ (.A0(_02207_),
    .A1(net1502),
    .S(_02220_),
    .X(_02227_));
 sky130_fd_sc_hd__clkbuf_1 _14844_ (.A(_02227_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _14845_ (.A0(_02209_),
    .A1(\cur_mb_mem[46][7] ),
    .S(_02220_),
    .X(_02228_));
 sky130_fd_sc_hd__clkbuf_1 _14846_ (.A(_02228_),
    .X(_00526_));
 sky130_fd_sc_hd__nand2_8 _14847_ (.A(_06259_),
    .B(_09319_),
    .Y(_02229_));
 sky130_fd_sc_hd__mux2_1 _14848_ (.A0(_02194_),
    .A1(net1120),
    .S(_02229_),
    .X(_02230_));
 sky130_fd_sc_hd__clkbuf_1 _14849_ (.A(_02230_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _14850_ (.A0(_02197_),
    .A1(\cur_mb_mem[47][1] ),
    .S(_02229_),
    .X(_02231_));
 sky130_fd_sc_hd__clkbuf_1 _14851_ (.A(_02231_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _14852_ (.A0(_02199_),
    .A1(net712),
    .S(_02229_),
    .X(_02232_));
 sky130_fd_sc_hd__clkbuf_1 _14853_ (.A(_02232_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _14854_ (.A0(_02201_),
    .A1(net1271),
    .S(_02229_),
    .X(_02233_));
 sky130_fd_sc_hd__clkbuf_1 _14855_ (.A(_02233_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _14856_ (.A0(_02203_),
    .A1(\cur_mb_mem[47][4] ),
    .S(_02229_),
    .X(_02234_));
 sky130_fd_sc_hd__clkbuf_1 _14857_ (.A(_02234_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _14858_ (.A0(_02205_),
    .A1(\cur_mb_mem[47][5] ),
    .S(_02229_),
    .X(_02235_));
 sky130_fd_sc_hd__clkbuf_1 _14859_ (.A(_02235_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _14860_ (.A0(_02207_),
    .A1(net1538),
    .S(_02229_),
    .X(_02236_));
 sky130_fd_sc_hd__clkbuf_1 _14861_ (.A(_02236_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _14862_ (.A0(_02209_),
    .A1(net1640),
    .S(_02229_),
    .X(_02237_));
 sky130_fd_sc_hd__clkbuf_1 _14863_ (.A(_02237_),
    .X(_00534_));
 sky130_fd_sc_hd__buf_4 _14864_ (.A(_05059_),
    .X(_02238_));
 sky130_fd_sc_hd__nand2_8 _14865_ (.A(_02238_),
    .B(_08883_),
    .Y(_02239_));
 sky130_fd_sc_hd__mux2_1 _14866_ (.A0(_02194_),
    .A1(net504),
    .S(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__clkbuf_1 _14867_ (.A(_02240_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _14868_ (.A0(_02197_),
    .A1(net835),
    .S(_02239_),
    .X(_02241_));
 sky130_fd_sc_hd__clkbuf_1 _14869_ (.A(_02241_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _14870_ (.A0(_02199_),
    .A1(net833),
    .S(_02239_),
    .X(_02242_));
 sky130_fd_sc_hd__clkbuf_1 _14871_ (.A(_02242_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _14872_ (.A0(_02201_),
    .A1(net711),
    .S(_02239_),
    .X(_02243_));
 sky130_fd_sc_hd__clkbuf_1 _14873_ (.A(_02243_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _14874_ (.A0(_02203_),
    .A1(net654),
    .S(_02239_),
    .X(_02244_));
 sky130_fd_sc_hd__clkbuf_1 _14875_ (.A(_02244_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _14876_ (.A0(_02205_),
    .A1(net618),
    .S(_02239_),
    .X(_02245_));
 sky130_fd_sc_hd__clkbuf_1 _14877_ (.A(_02245_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _14878_ (.A0(_02207_),
    .A1(net1419),
    .S(_02239_),
    .X(_02246_));
 sky130_fd_sc_hd__clkbuf_1 _14879_ (.A(_02246_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _14880_ (.A0(_02209_),
    .A1(net1199),
    .S(_02239_),
    .X(_02247_));
 sky130_fd_sc_hd__clkbuf_1 _14881_ (.A(_02247_),
    .X(_00542_));
 sky130_fd_sc_hd__nand3_4 _14882_ (.A(_02238_),
    .B(_05994_),
    .C(_08979_),
    .Y(_02248_));
 sky130_fd_sc_hd__mux2_1 _14883_ (.A0(_02194_),
    .A1(net495),
    .S(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__clkbuf_1 _14884_ (.A(_02249_),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _14885_ (.A0(_02197_),
    .A1(net649),
    .S(_02248_),
    .X(_02250_));
 sky130_fd_sc_hd__clkbuf_1 _14886_ (.A(_02250_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _14887_ (.A0(_02199_),
    .A1(net752),
    .S(_02248_),
    .X(_02251_));
 sky130_fd_sc_hd__clkbuf_1 _14888_ (.A(_02251_),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _14889_ (.A0(_02201_),
    .A1(net772),
    .S(_02248_),
    .X(_02252_));
 sky130_fd_sc_hd__clkbuf_1 _14890_ (.A(_02252_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _14891_ (.A0(_02203_),
    .A1(net634),
    .S(_02248_),
    .X(_02253_));
 sky130_fd_sc_hd__clkbuf_1 _14892_ (.A(_02253_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _14893_ (.A0(_02205_),
    .A1(net713),
    .S(_02248_),
    .X(_02254_));
 sky130_fd_sc_hd__clkbuf_1 _14894_ (.A(_02254_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _14895_ (.A0(_02207_),
    .A1(net1295),
    .S(_02248_),
    .X(_02255_));
 sky130_fd_sc_hd__clkbuf_1 _14896_ (.A(_02255_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _14897_ (.A0(_02209_),
    .A1(net1329),
    .S(_02248_),
    .X(_02256_));
 sky130_fd_sc_hd__clkbuf_1 _14898_ (.A(_02256_),
    .X(_00550_));
 sky130_fd_sc_hd__nand2_8 _14899_ (.A(_06172_),
    .B(_09319_),
    .Y(_02257_));
 sky130_fd_sc_hd__mux2_1 _14900_ (.A0(_02194_),
    .A1(net1611),
    .S(_02257_),
    .X(_02258_));
 sky130_fd_sc_hd__clkbuf_1 _14901_ (.A(_02258_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _14902_ (.A0(_02197_),
    .A1(net542),
    .S(_02257_),
    .X(_02259_));
 sky130_fd_sc_hd__clkbuf_1 _14903_ (.A(_02259_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _14904_ (.A0(_02199_),
    .A1(net1595),
    .S(_02257_),
    .X(_02260_));
 sky130_fd_sc_hd__clkbuf_1 _14905_ (.A(_02260_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _14906_ (.A0(_02201_),
    .A1(net1146),
    .S(_02257_),
    .X(_02261_));
 sky130_fd_sc_hd__clkbuf_1 _14907_ (.A(_02261_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _14908_ (.A0(_02203_),
    .A1(net1683),
    .S(_02257_),
    .X(_02262_));
 sky130_fd_sc_hd__clkbuf_1 _14909_ (.A(_02262_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _14910_ (.A0(_02205_),
    .A1(net1705),
    .S(_02257_),
    .X(_02263_));
 sky130_fd_sc_hd__clkbuf_1 _14911_ (.A(_02263_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _14912_ (.A0(_02207_),
    .A1(net1790),
    .S(_02257_),
    .X(_02264_));
 sky130_fd_sc_hd__clkbuf_1 _14913_ (.A(_02264_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _14914_ (.A0(_02209_),
    .A1(net1210),
    .S(_02257_),
    .X(_02265_));
 sky130_fd_sc_hd__clkbuf_1 _14915_ (.A(_02265_),
    .X(_00558_));
 sky130_fd_sc_hd__buf_8 _14916_ (.A(_06064_),
    .X(_02266_));
 sky130_fd_sc_hd__and3_1 _14917_ (.A(_02238_),
    .B(_02266_),
    .C(_09037_),
    .X(_02267_));
 sky130_fd_sc_hd__buf_6 _14918_ (.A(_02267_),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _14919_ (.A0(net1298),
    .A1(_08531_),
    .S(_02268_),
    .X(_02269_));
 sky130_fd_sc_hd__clkbuf_1 _14920_ (.A(_02269_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _14921_ (.A0(net1039),
    .A1(_08536_),
    .S(_02268_),
    .X(_02270_));
 sky130_fd_sc_hd__clkbuf_1 _14922_ (.A(_02270_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _14923_ (.A0(\cur_mb_mem[51][2] ),
    .A1(_08539_),
    .S(_02268_),
    .X(_02271_));
 sky130_fd_sc_hd__clkbuf_1 _14924_ (.A(_02271_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _14925_ (.A0(net678),
    .A1(_08542_),
    .S(_02268_),
    .X(_02272_));
 sky130_fd_sc_hd__clkbuf_1 _14926_ (.A(_02272_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _14927_ (.A0(net1294),
    .A1(_08545_),
    .S(_02268_),
    .X(_02273_));
 sky130_fd_sc_hd__clkbuf_1 _14928_ (.A(_02273_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _14929_ (.A0(net1038),
    .A1(_08548_),
    .S(_02268_),
    .X(_02274_));
 sky130_fd_sc_hd__clkbuf_1 _14930_ (.A(_02274_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _14931_ (.A0(net1263),
    .A1(_08551_),
    .S(_02268_),
    .X(_02275_));
 sky130_fd_sc_hd__clkbuf_1 _14932_ (.A(_02275_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _14933_ (.A0(net1963),
    .A1(_08554_),
    .S(_02268_),
    .X(_02276_));
 sky130_fd_sc_hd__clkbuf_1 _14934_ (.A(_02276_),
    .X(_00566_));
 sky130_fd_sc_hd__nand2_8 _14935_ (.A(_06241_),
    .B(_09319_),
    .Y(_02277_));
 sky130_fd_sc_hd__mux2_1 _14936_ (.A0(_02194_),
    .A1(net1487),
    .S(_02277_),
    .X(_02278_));
 sky130_fd_sc_hd__clkbuf_1 _14937_ (.A(_02278_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _14938_ (.A0(_02197_),
    .A1(net675),
    .S(_02277_),
    .X(_02279_));
 sky130_fd_sc_hd__clkbuf_1 _14939_ (.A(_02279_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _14940_ (.A0(_02199_),
    .A1(net1190),
    .S(_02277_),
    .X(_02280_));
 sky130_fd_sc_hd__clkbuf_1 _14941_ (.A(_02280_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _14942_ (.A0(_02201_),
    .A1(net1282),
    .S(_02277_),
    .X(_02281_));
 sky130_fd_sc_hd__clkbuf_1 _14943_ (.A(_02281_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _14944_ (.A0(_02203_),
    .A1(net1065),
    .S(_02277_),
    .X(_02282_));
 sky130_fd_sc_hd__clkbuf_1 _14945_ (.A(_02282_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _14946_ (.A0(_02205_),
    .A1(net787),
    .S(_02277_),
    .X(_02283_));
 sky130_fd_sc_hd__clkbuf_1 _14947_ (.A(_02283_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _14948_ (.A0(_02207_),
    .A1(net1782),
    .S(_02277_),
    .X(_02284_));
 sky130_fd_sc_hd__clkbuf_1 _14949_ (.A(_02284_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _14950_ (.A0(_02209_),
    .A1(net1546),
    .S(_02277_),
    .X(_02285_));
 sky130_fd_sc_hd__clkbuf_1 _14951_ (.A(_02285_),
    .X(_00574_));
 sky130_fd_sc_hd__buf_8 _14952_ (.A(_06133_),
    .X(_02286_));
 sky130_fd_sc_hd__and3_1 _14953_ (.A(_02238_),
    .B(_02286_),
    .C(_09037_),
    .X(_02287_));
 sky130_fd_sc_hd__buf_8 _14954_ (.A(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _14955_ (.A0(net1083),
    .A1(_08531_),
    .S(_02288_),
    .X(_02289_));
 sky130_fd_sc_hd__clkbuf_1 _14956_ (.A(_02289_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _14957_ (.A0(net463),
    .A1(_08536_),
    .S(_02288_),
    .X(_02290_));
 sky130_fd_sc_hd__clkbuf_1 _14958_ (.A(_02290_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _14959_ (.A0(net928),
    .A1(_08539_),
    .S(_02288_),
    .X(_02291_));
 sky130_fd_sc_hd__clkbuf_1 _14960_ (.A(_02291_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _14961_ (.A0(net1211),
    .A1(_08542_),
    .S(_02288_),
    .X(_02292_));
 sky130_fd_sc_hd__clkbuf_1 _14962_ (.A(_02292_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _14963_ (.A0(net1723),
    .A1(_08545_),
    .S(_02288_),
    .X(_02293_));
 sky130_fd_sc_hd__clkbuf_1 _14964_ (.A(_02293_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _14965_ (.A0(net1012),
    .A1(_08548_),
    .S(_02288_),
    .X(_02294_));
 sky130_fd_sc_hd__clkbuf_1 _14966_ (.A(_02294_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _14967_ (.A0(net1729),
    .A1(_08551_),
    .S(_02288_),
    .X(_02295_));
 sky130_fd_sc_hd__clkbuf_1 _14968_ (.A(_02295_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _14969_ (.A0(net999),
    .A1(_08554_),
    .S(_02288_),
    .X(_02296_));
 sky130_fd_sc_hd__clkbuf_1 _14970_ (.A(_02296_),
    .X(_00582_));
 sky130_fd_sc_hd__buf_6 _14971_ (.A(_06187_),
    .X(_02297_));
 sky130_fd_sc_hd__and3_1 _14972_ (.A(_02238_),
    .B(_02297_),
    .C(_09037_),
    .X(_02298_));
 sky130_fd_sc_hd__buf_6 _14973_ (.A(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__mux2_1 _14974_ (.A0(net1694),
    .A1(_08531_),
    .S(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__clkbuf_1 _14975_ (.A(_02300_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _14976_ (.A0(net348),
    .A1(_08536_),
    .S(_02299_),
    .X(_02301_));
 sky130_fd_sc_hd__clkbuf_1 _14977_ (.A(_02301_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _14978_ (.A0(net1976),
    .A1(_08539_),
    .S(_02299_),
    .X(_02302_));
 sky130_fd_sc_hd__clkbuf_1 _14979_ (.A(_02302_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _14980_ (.A0(net714),
    .A1(_08542_),
    .S(_02299_),
    .X(_02303_));
 sky130_fd_sc_hd__clkbuf_1 _14981_ (.A(_02303_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _14982_ (.A0(net625),
    .A1(_08545_),
    .S(_02299_),
    .X(_02304_));
 sky130_fd_sc_hd__clkbuf_1 _14983_ (.A(_02304_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _14984_ (.A0(net530),
    .A1(_08548_),
    .S(_02299_),
    .X(_02305_));
 sky130_fd_sc_hd__clkbuf_1 _14985_ (.A(_02305_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _14986_ (.A0(net1972),
    .A1(_08551_),
    .S(_02299_),
    .X(_02306_));
 sky130_fd_sc_hd__clkbuf_1 _14987_ (.A(_02306_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _14988_ (.A0(net551),
    .A1(_08554_),
    .S(_02299_),
    .X(_02307_));
 sky130_fd_sc_hd__clkbuf_1 _14989_ (.A(_02307_),
    .X(_00590_));
 sky130_fd_sc_hd__and3_1 _14990_ (.A(_02238_),
    .B(_08839_),
    .C(_09037_),
    .X(_02308_));
 sky130_fd_sc_hd__buf_6 _14991_ (.A(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _14992_ (.A0(net696),
    .A1(_08531_),
    .S(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__clkbuf_1 _14993_ (.A(_02310_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _14994_ (.A0(net423),
    .A1(_08536_),
    .S(_02309_),
    .X(_02311_));
 sky130_fd_sc_hd__clkbuf_1 _14995_ (.A(_02311_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _14996_ (.A0(net446),
    .A1(_08539_),
    .S(_02309_),
    .X(_02312_));
 sky130_fd_sc_hd__clkbuf_1 _14997_ (.A(_02312_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _14998_ (.A0(net815),
    .A1(_08542_),
    .S(_02309_),
    .X(_02313_));
 sky130_fd_sc_hd__clkbuf_1 _14999_ (.A(_02313_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _15000_ (.A0(net1157),
    .A1(_08545_),
    .S(_02309_),
    .X(_02314_));
 sky130_fd_sc_hd__clkbuf_1 _15001_ (.A(_02314_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _15002_ (.A0(net1266),
    .A1(_08548_),
    .S(_02309_),
    .X(_02315_));
 sky130_fd_sc_hd__clkbuf_1 _15003_ (.A(_02315_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _15004_ (.A0(net624),
    .A1(_08551_),
    .S(_02309_),
    .X(_02316_));
 sky130_fd_sc_hd__clkbuf_1 _15005_ (.A(_02316_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _15006_ (.A0(net967),
    .A1(_08554_),
    .S(_02309_),
    .X(_02317_));
 sky130_fd_sc_hd__clkbuf_1 _15007_ (.A(_02317_),
    .X(_00598_));
 sky130_fd_sc_hd__nand2_8 _15008_ (.A(_06351_),
    .B(_09319_),
    .Y(_02318_));
 sky130_fd_sc_hd__mux2_1 _15009_ (.A0(_02194_),
    .A1(net1258),
    .S(_02318_),
    .X(_02319_));
 sky130_fd_sc_hd__clkbuf_1 _15010_ (.A(_02319_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _15011_ (.A0(_02197_),
    .A1(net955),
    .S(_02318_),
    .X(_02320_));
 sky130_fd_sc_hd__clkbuf_1 _15012_ (.A(_02320_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _15013_ (.A0(_02199_),
    .A1(net1352),
    .S(_02318_),
    .X(_02321_));
 sky130_fd_sc_hd__clkbuf_1 _15014_ (.A(_02321_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _15015_ (.A0(_02201_),
    .A1(net1501),
    .S(_02318_),
    .X(_02322_));
 sky130_fd_sc_hd__clkbuf_1 _15016_ (.A(_02322_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _15017_ (.A0(_02203_),
    .A1(net840),
    .S(_02318_),
    .X(_02323_));
 sky130_fd_sc_hd__clkbuf_1 _15018_ (.A(_02323_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _15019_ (.A0(_02205_),
    .A1(net707),
    .S(_02318_),
    .X(_02324_));
 sky130_fd_sc_hd__clkbuf_1 _15020_ (.A(_02324_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _15021_ (.A0(_02207_),
    .A1(net1759),
    .S(_02318_),
    .X(_02325_));
 sky130_fd_sc_hd__clkbuf_1 _15022_ (.A(_02325_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _15023_ (.A0(_02209_),
    .A1(\cur_mb_mem[56][7] ),
    .S(_02318_),
    .X(_02326_));
 sky130_fd_sc_hd__clkbuf_1 _15024_ (.A(_02326_),
    .X(_00606_));
 sky130_fd_sc_hd__clkbuf_8 _15025_ (.A(net97),
    .X(_02327_));
 sky130_fd_sc_hd__buf_12 _15026_ (.A(_02327_),
    .X(_02328_));
 sky130_fd_sc_hd__and3_1 _15027_ (.A(_02238_),
    .B(_05912_),
    .C(_09037_),
    .X(_02329_));
 sky130_fd_sc_hd__buf_8 _15028_ (.A(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__mux2_1 _15029_ (.A0(net320),
    .A1(_02328_),
    .S(_02330_),
    .X(_02331_));
 sky130_fd_sc_hd__clkbuf_1 _15030_ (.A(_02331_),
    .X(_00607_));
 sky130_fd_sc_hd__buf_4 _15031_ (.A(net98),
    .X(_02332_));
 sky130_fd_sc_hd__buf_8 _15032_ (.A(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__mux2_1 _15033_ (.A0(net385),
    .A1(_02333_),
    .S(_02330_),
    .X(_02334_));
 sky130_fd_sc_hd__clkbuf_1 _15034_ (.A(_02334_),
    .X(_00608_));
 sky130_fd_sc_hd__clkbuf_8 _15035_ (.A(net99),
    .X(_02335_));
 sky130_fd_sc_hd__clkbuf_16 _15036_ (.A(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__mux2_1 _15037_ (.A0(net1627),
    .A1(_02336_),
    .S(_02330_),
    .X(_02337_));
 sky130_fd_sc_hd__clkbuf_1 _15038_ (.A(_02337_),
    .X(_00609_));
 sky130_fd_sc_hd__clkbuf_8 _15039_ (.A(net100),
    .X(_02338_));
 sky130_fd_sc_hd__clkbuf_16 _15040_ (.A(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__mux2_1 _15041_ (.A0(net407),
    .A1(_02339_),
    .S(_02330_),
    .X(_02340_));
 sky130_fd_sc_hd__clkbuf_1 _15042_ (.A(_02340_),
    .X(_00610_));
 sky130_fd_sc_hd__buf_8 _15043_ (.A(net101),
    .X(_02341_));
 sky130_fd_sc_hd__clkbuf_16 _15044_ (.A(_02341_),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _15045_ (.A0(net393),
    .A1(_02342_),
    .S(_02330_),
    .X(_02343_));
 sky130_fd_sc_hd__clkbuf_1 _15046_ (.A(_02343_),
    .X(_00611_));
 sky130_fd_sc_hd__buf_8 _15047_ (.A(net102),
    .X(_02344_));
 sky130_fd_sc_hd__clkbuf_16 _15048_ (.A(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__mux2_1 _15049_ (.A0(net642),
    .A1(_02345_),
    .S(_02330_),
    .X(_02346_));
 sky130_fd_sc_hd__clkbuf_1 _15050_ (.A(_02346_),
    .X(_00612_));
 sky130_fd_sc_hd__clkbuf_8 _15051_ (.A(net103),
    .X(_02347_));
 sky130_fd_sc_hd__buf_6 _15052_ (.A(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__mux2_1 _15053_ (.A0(net1072),
    .A1(_02348_),
    .S(_02330_),
    .X(_02349_));
 sky130_fd_sc_hd__clkbuf_1 _15054_ (.A(_02349_),
    .X(_00613_));
 sky130_fd_sc_hd__buf_4 _15055_ (.A(net104),
    .X(_02350_));
 sky130_fd_sc_hd__clkbuf_8 _15056_ (.A(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__mux2_1 _15057_ (.A0(net761),
    .A1(_02351_),
    .S(_02330_),
    .X(_02352_));
 sky130_fd_sc_hd__clkbuf_1 _15058_ (.A(_02352_),
    .X(_00614_));
 sky130_fd_sc_hd__buf_8 _15059_ (.A(_06035_),
    .X(_02353_));
 sky130_fd_sc_hd__and3_1 _15060_ (.A(_02238_),
    .B(_02353_),
    .C(_09037_),
    .X(_02354_));
 sky130_fd_sc_hd__buf_8 _15061_ (.A(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__mux2_1 _15062_ (.A0(net416),
    .A1(_02328_),
    .S(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__clkbuf_1 _15063_ (.A(_02356_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _15064_ (.A0(net331),
    .A1(_02333_),
    .S(_02355_),
    .X(_02357_));
 sky130_fd_sc_hd__clkbuf_1 _15065_ (.A(_02357_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _15066_ (.A0(net938),
    .A1(_02336_),
    .S(_02355_),
    .X(_02358_));
 sky130_fd_sc_hd__clkbuf_1 _15067_ (.A(_02358_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _15068_ (.A0(net461),
    .A1(_02339_),
    .S(_02355_),
    .X(_02359_));
 sky130_fd_sc_hd__clkbuf_1 _15069_ (.A(_02359_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _15070_ (.A0(net522),
    .A1(_02342_),
    .S(_02355_),
    .X(_02360_));
 sky130_fd_sc_hd__clkbuf_1 _15071_ (.A(_02360_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _15072_ (.A0(net429),
    .A1(_02345_),
    .S(_02355_),
    .X(_02361_));
 sky130_fd_sc_hd__clkbuf_1 _15073_ (.A(_02361_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _15074_ (.A0(net1020),
    .A1(_02348_),
    .S(_02355_),
    .X(_02362_));
 sky130_fd_sc_hd__clkbuf_1 _15075_ (.A(_02362_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _15076_ (.A0(net1050),
    .A1(_02351_),
    .S(_02355_),
    .X(_02363_));
 sky130_fd_sc_hd__clkbuf_1 _15077_ (.A(_02363_),
    .X(_00622_));
 sky130_fd_sc_hd__and3_1 _15078_ (.A(_02238_),
    .B(_06049_),
    .C(_09037_),
    .X(_02364_));
 sky130_fd_sc_hd__buf_4 _15079_ (.A(_02364_),
    .X(_02365_));
 sky130_fd_sc_hd__mux2_1 _15080_ (.A0(net561),
    .A1(_02328_),
    .S(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__clkbuf_1 _15081_ (.A(_02366_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _15082_ (.A0(net377),
    .A1(_02333_),
    .S(_02365_),
    .X(_02367_));
 sky130_fd_sc_hd__clkbuf_1 _15083_ (.A(_02367_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _15084_ (.A0(net524),
    .A1(_02336_),
    .S(_02365_),
    .X(_02368_));
 sky130_fd_sc_hd__clkbuf_1 _15085_ (.A(_02368_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _15086_ (.A0(net560),
    .A1(_02339_),
    .S(_02365_),
    .X(_02369_));
 sky130_fd_sc_hd__clkbuf_1 _15087_ (.A(_02369_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _15088_ (.A0(net656),
    .A1(_02342_),
    .S(_02365_),
    .X(_02370_));
 sky130_fd_sc_hd__clkbuf_1 _15089_ (.A(_02370_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _15090_ (.A0(net896),
    .A1(_02345_),
    .S(_02365_),
    .X(_02371_));
 sky130_fd_sc_hd__clkbuf_1 _15091_ (.A(_02371_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _15092_ (.A0(net600),
    .A1(_02348_),
    .S(_02365_),
    .X(_02372_));
 sky130_fd_sc_hd__clkbuf_1 _15093_ (.A(_02372_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _15094_ (.A0(net1625),
    .A1(_02351_),
    .S(_02365_),
    .X(_02373_));
 sky130_fd_sc_hd__clkbuf_1 _15095_ (.A(_02373_),
    .X(_00630_));
 sky130_fd_sc_hd__buf_8 _15096_ (.A(_05989_),
    .X(_02374_));
 sky130_fd_sc_hd__and3_1 _15097_ (.A(_02238_),
    .B(_02374_),
    .C(_09037_),
    .X(_02375_));
 sky130_fd_sc_hd__clkbuf_16 _15098_ (.A(_02375_),
    .X(_02376_));
 sky130_fd_sc_hd__mux2_1 _15099_ (.A0(net577),
    .A1(_02328_),
    .S(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__clkbuf_1 _15100_ (.A(_02377_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _15101_ (.A0(net610),
    .A1(_02333_),
    .S(_02376_),
    .X(_02378_));
 sky130_fd_sc_hd__clkbuf_1 _15102_ (.A(_02378_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _15103_ (.A0(net408),
    .A1(_02336_),
    .S(_02376_),
    .X(_02379_));
 sky130_fd_sc_hd__clkbuf_1 _15104_ (.A(_02379_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _15105_ (.A0(net343),
    .A1(_02339_),
    .S(_02376_),
    .X(_02380_));
 sky130_fd_sc_hd__clkbuf_1 _15106_ (.A(_02380_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _15107_ (.A0(net471),
    .A1(_02342_),
    .S(_02376_),
    .X(_02381_));
 sky130_fd_sc_hd__clkbuf_1 _15108_ (.A(_02381_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _15109_ (.A0(net1031),
    .A1(_02345_),
    .S(_02376_),
    .X(_02382_));
 sky130_fd_sc_hd__clkbuf_1 _15110_ (.A(_02382_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _15111_ (.A0(net1064),
    .A1(_02348_),
    .S(_02376_),
    .X(_02383_));
 sky130_fd_sc_hd__clkbuf_1 _15112_ (.A(_02383_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _15113_ (.A0(net791),
    .A1(_02351_),
    .S(_02376_),
    .X(_02384_));
 sky130_fd_sc_hd__clkbuf_1 _15114_ (.A(_02384_),
    .X(_00638_));
 sky130_fd_sc_hd__and3_1 _15115_ (.A(_05059_),
    .B(_09025_),
    .C(_09037_),
    .X(_02385_));
 sky130_fd_sc_hd__buf_8 _15116_ (.A(_02385_),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _15117_ (.A0(\cur_mb_mem[61][0] ),
    .A1(_02328_),
    .S(_02386_),
    .X(_02387_));
 sky130_fd_sc_hd__clkbuf_1 _15118_ (.A(_02387_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _15119_ (.A0(net1310),
    .A1(_02333_),
    .S(_02386_),
    .X(_02388_));
 sky130_fd_sc_hd__clkbuf_1 _15120_ (.A(_02388_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _15121_ (.A0(net1139),
    .A1(_02336_),
    .S(_02386_),
    .X(_02389_));
 sky130_fd_sc_hd__clkbuf_1 _15122_ (.A(_02389_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _15123_ (.A0(net1385),
    .A1(_02339_),
    .S(_02386_),
    .X(_02390_));
 sky130_fd_sc_hd__clkbuf_1 _15124_ (.A(_02390_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _15125_ (.A0(net1121),
    .A1(_02342_),
    .S(_02386_),
    .X(_02391_));
 sky130_fd_sc_hd__clkbuf_1 _15126_ (.A(_02391_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _15127_ (.A0(net994),
    .A1(_02345_),
    .S(_02386_),
    .X(_02392_));
 sky130_fd_sc_hd__clkbuf_1 _15128_ (.A(_02392_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _15129_ (.A0(net943),
    .A1(_02348_),
    .S(_02386_),
    .X(_02393_));
 sky130_fd_sc_hd__clkbuf_1 _15130_ (.A(_02393_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _15131_ (.A0(net1005),
    .A1(_02351_),
    .S(_02386_),
    .X(_02394_));
 sky130_fd_sc_hd__clkbuf_1 _15132_ (.A(_02394_),
    .X(_00646_));
 sky130_fd_sc_hd__buf_2 _15133_ (.A(_08900_),
    .X(_02395_));
 sky130_fd_sc_hd__and3_1 _15134_ (.A(_05059_),
    .B(_09036_),
    .C(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__buf_6 _15135_ (.A(_02396_),
    .X(_02397_));
 sky130_fd_sc_hd__mux2_1 _15136_ (.A0(net648),
    .A1(_02328_),
    .S(_02397_),
    .X(_02398_));
 sky130_fd_sc_hd__clkbuf_1 _15137_ (.A(_02398_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _15138_ (.A0(net1391),
    .A1(_02333_),
    .S(_02397_),
    .X(_02399_));
 sky130_fd_sc_hd__clkbuf_1 _15139_ (.A(_02399_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _15140_ (.A0(net518),
    .A1(_02336_),
    .S(_02397_),
    .X(_02400_));
 sky130_fd_sc_hd__clkbuf_1 _15141_ (.A(_02400_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _15142_ (.A0(net684),
    .A1(_02339_),
    .S(_02397_),
    .X(_02401_));
 sky130_fd_sc_hd__clkbuf_1 _15143_ (.A(_02401_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _15144_ (.A0(net812),
    .A1(_02342_),
    .S(_02397_),
    .X(_02402_));
 sky130_fd_sc_hd__clkbuf_1 _15145_ (.A(_02402_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _15146_ (.A0(net563),
    .A1(_02345_),
    .S(_02397_),
    .X(_02403_));
 sky130_fd_sc_hd__clkbuf_1 _15147_ (.A(_02403_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _15148_ (.A0(net864),
    .A1(_02348_),
    .S(_02397_),
    .X(_02404_));
 sky130_fd_sc_hd__clkbuf_1 _15149_ (.A(_02404_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _15150_ (.A0(net1117),
    .A1(_02351_),
    .S(_02397_),
    .X(_02405_));
 sky130_fd_sc_hd__clkbuf_1 _15151_ (.A(_02405_),
    .X(_00654_));
 sky130_fd_sc_hd__clkbuf_8 _15152_ (.A(_04424_),
    .X(_02406_));
 sky130_fd_sc_hd__and3_1 _15153_ (.A(_02406_),
    .B(_05059_),
    .C(_02395_),
    .X(_02407_));
 sky130_fd_sc_hd__buf_4 _15154_ (.A(_02407_),
    .X(_02408_));
 sky130_fd_sc_hd__mux2_1 _15155_ (.A0(net438),
    .A1(_02328_),
    .S(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__clkbuf_1 _15156_ (.A(_02409_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _15157_ (.A0(net783),
    .A1(_02333_),
    .S(_02408_),
    .X(_02410_));
 sky130_fd_sc_hd__clkbuf_1 _15158_ (.A(_02410_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _15159_ (.A0(net397),
    .A1(_02336_),
    .S(_02408_),
    .X(_02411_));
 sky130_fd_sc_hd__clkbuf_1 _15160_ (.A(_02411_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _15161_ (.A0(net411),
    .A1(_02339_),
    .S(_02408_),
    .X(_02412_));
 sky130_fd_sc_hd__clkbuf_1 _15162_ (.A(_02412_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _15163_ (.A0(net669),
    .A1(_02342_),
    .S(_02408_),
    .X(_02413_));
 sky130_fd_sc_hd__clkbuf_1 _15164_ (.A(_02413_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _15165_ (.A0(net442),
    .A1(_02345_),
    .S(_02408_),
    .X(_02414_));
 sky130_fd_sc_hd__clkbuf_1 _15166_ (.A(_02414_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _15167_ (.A0(net1006),
    .A1(_02348_),
    .S(_02408_),
    .X(_02415_));
 sky130_fd_sc_hd__clkbuf_1 _15168_ (.A(_02415_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _15169_ (.A0(net1178),
    .A1(_02351_),
    .S(_02408_),
    .X(_02416_));
 sky130_fd_sc_hd__clkbuf_1 _15170_ (.A(_02416_),
    .X(_00662_));
 sky130_fd_sc_hd__nand2_8 _15171_ (.A(_06024_),
    .B(_08883_),
    .Y(_02417_));
 sky130_fd_sc_hd__mux2_1 _15172_ (.A0(_02194_),
    .A1(net904),
    .S(_02417_),
    .X(_02418_));
 sky130_fd_sc_hd__clkbuf_1 _15173_ (.A(_02418_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _15174_ (.A0(_02197_),
    .A1(net483),
    .S(_02417_),
    .X(_02419_));
 sky130_fd_sc_hd__clkbuf_1 _15175_ (.A(_02419_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _15176_ (.A0(_02199_),
    .A1(net1098),
    .S(_02417_),
    .X(_02420_));
 sky130_fd_sc_hd__clkbuf_1 _15177_ (.A(_02420_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _15178_ (.A0(_02201_),
    .A1(net683),
    .S(_02417_),
    .X(_02421_));
 sky130_fd_sc_hd__clkbuf_1 _15179_ (.A(_02421_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _15180_ (.A0(_02203_),
    .A1(net736),
    .S(_02417_),
    .X(_02422_));
 sky130_fd_sc_hd__clkbuf_1 _15181_ (.A(_02422_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _15182_ (.A0(_02205_),
    .A1(net1116),
    .S(_02417_),
    .X(_02423_));
 sky130_fd_sc_hd__clkbuf_1 _15183_ (.A(_02423_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _15184_ (.A0(_02207_),
    .A1(\cur_mb_mem[64][6] ),
    .S(_02417_),
    .X(_02424_));
 sky130_fd_sc_hd__clkbuf_1 _15185_ (.A(_02424_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _15186_ (.A0(_02209_),
    .A1(net1442),
    .S(_02417_),
    .X(_02425_));
 sky130_fd_sc_hd__clkbuf_1 _15187_ (.A(_02425_),
    .X(_00670_));
 sky130_fd_sc_hd__clkbuf_4 _15188_ (.A(_09132_),
    .X(_02426_));
 sky130_fd_sc_hd__nand2_8 _15189_ (.A(_06483_),
    .B(_09319_),
    .Y(_02427_));
 sky130_fd_sc_hd__mux2_1 _15190_ (.A0(_02426_),
    .A1(net1060),
    .S(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__clkbuf_1 _15191_ (.A(_02428_),
    .X(_00671_));
 sky130_fd_sc_hd__buf_4 _15192_ (.A(_09136_),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _15193_ (.A0(_02429_),
    .A1(\cur_mb_mem[65][1] ),
    .S(_02427_),
    .X(_02430_));
 sky130_fd_sc_hd__clkbuf_1 _15194_ (.A(_02430_),
    .X(_00672_));
 sky130_fd_sc_hd__buf_4 _15195_ (.A(_09139_),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _15196_ (.A0(_02431_),
    .A1(net1482),
    .S(_02427_),
    .X(_02432_));
 sky130_fd_sc_hd__clkbuf_1 _15197_ (.A(_02432_),
    .X(_00673_));
 sky130_fd_sc_hd__clkbuf_4 _15198_ (.A(_09142_),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_1 _15199_ (.A0(_02433_),
    .A1(net1055),
    .S(_02427_),
    .X(_02434_));
 sky130_fd_sc_hd__clkbuf_1 _15200_ (.A(_02434_),
    .X(_00674_));
 sky130_fd_sc_hd__clkbuf_4 _15201_ (.A(_09145_),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _15202_ (.A0(_02435_),
    .A1(net1674),
    .S(_02427_),
    .X(_02436_));
 sky130_fd_sc_hd__clkbuf_1 _15203_ (.A(_02436_),
    .X(_00675_));
 sky130_fd_sc_hd__clkbuf_4 _15204_ (.A(_09148_),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _15205_ (.A0(_02437_),
    .A1(net1696),
    .S(_02427_),
    .X(_02438_));
 sky130_fd_sc_hd__clkbuf_1 _15206_ (.A(_02438_),
    .X(_00676_));
 sky130_fd_sc_hd__clkbuf_4 _15207_ (.A(_09151_),
    .X(_02439_));
 sky130_fd_sc_hd__mux2_1 _15208_ (.A0(_02439_),
    .A1(net1806),
    .S(_02427_),
    .X(_02440_));
 sky130_fd_sc_hd__clkbuf_1 _15209_ (.A(_02440_),
    .X(_00677_));
 sky130_fd_sc_hd__buf_4 _15210_ (.A(_09154_),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _15211_ (.A0(_02441_),
    .A1(\cur_mb_mem[65][7] ),
    .S(_02427_),
    .X(_02442_));
 sky130_fd_sc_hd__clkbuf_1 _15212_ (.A(_02442_),
    .X(_00678_));
 sky130_fd_sc_hd__buf_12 _15213_ (.A(_08958_),
    .X(_02443_));
 sky130_fd_sc_hd__nand2_8 _15214_ (.A(_06368_),
    .B(_02443_),
    .Y(_02444_));
 sky130_fd_sc_hd__mux2_1 _15215_ (.A0(_02426_),
    .A1(net1733),
    .S(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__clkbuf_1 _15216_ (.A(_02445_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _15217_ (.A0(_02429_),
    .A1(net1378),
    .S(_02444_),
    .X(_02446_));
 sky130_fd_sc_hd__clkbuf_1 _15218_ (.A(_02446_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _15219_ (.A0(_02431_),
    .A1(net1425),
    .S(_02444_),
    .X(_02447_));
 sky130_fd_sc_hd__clkbuf_1 _15220_ (.A(_02447_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _15221_ (.A0(_02433_),
    .A1(net1280),
    .S(_02444_),
    .X(_02448_));
 sky130_fd_sc_hd__clkbuf_1 _15222_ (.A(_02448_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _15223_ (.A0(_02435_),
    .A1(net1369),
    .S(_02444_),
    .X(_02449_));
 sky130_fd_sc_hd__clkbuf_1 _15224_ (.A(_02449_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _15225_ (.A0(_02437_),
    .A1(net1220),
    .S(_02444_),
    .X(_02450_));
 sky130_fd_sc_hd__clkbuf_1 _15226_ (.A(_02450_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _15227_ (.A0(_02439_),
    .A1(net1003),
    .S(_02444_),
    .X(_02451_));
 sky130_fd_sc_hd__clkbuf_1 _15228_ (.A(_02451_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _15229_ (.A0(_02441_),
    .A1(net1243),
    .S(_02444_),
    .X(_02452_));
 sky130_fd_sc_hd__clkbuf_1 _15230_ (.A(_02452_),
    .X(_00686_));
 sky130_fd_sc_hd__nand2_8 _15231_ (.A(_06429_),
    .B(_02443_),
    .Y(_02453_));
 sky130_fd_sc_hd__mux2_1 _15232_ (.A0(_02426_),
    .A1(\cur_mb_mem[67][0] ),
    .S(_02453_),
    .X(_02454_));
 sky130_fd_sc_hd__clkbuf_1 _15233_ (.A(_02454_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _15234_ (.A0(_02429_),
    .A1(net982),
    .S(_02453_),
    .X(_02455_));
 sky130_fd_sc_hd__clkbuf_1 _15235_ (.A(_02455_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _15236_ (.A0(_02431_),
    .A1(\cur_mb_mem[67][2] ),
    .S(_02453_),
    .X(_02456_));
 sky130_fd_sc_hd__clkbuf_1 _15237_ (.A(_02456_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _15238_ (.A0(_02433_),
    .A1(\cur_mb_mem[67][3] ),
    .S(_02453_),
    .X(_02457_));
 sky130_fd_sc_hd__clkbuf_1 _15239_ (.A(_02457_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _15240_ (.A0(_02435_),
    .A1(net1776),
    .S(_02453_),
    .X(_02458_));
 sky130_fd_sc_hd__clkbuf_1 _15241_ (.A(_02458_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _15242_ (.A0(_02437_),
    .A1(net1554),
    .S(_02453_),
    .X(_02459_));
 sky130_fd_sc_hd__clkbuf_1 _15243_ (.A(_02459_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _15244_ (.A0(_02439_),
    .A1(net1567),
    .S(_02453_),
    .X(_02460_));
 sky130_fd_sc_hd__clkbuf_1 _15245_ (.A(_02460_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _15246_ (.A0(_02441_),
    .A1(\cur_mb_mem[67][7] ),
    .S(_02453_),
    .X(_02461_));
 sky130_fd_sc_hd__clkbuf_1 _15247_ (.A(_02461_),
    .X(_00694_));
 sky130_fd_sc_hd__nand2_8 _15248_ (.A(_06234_),
    .B(_02443_),
    .Y(_02462_));
 sky130_fd_sc_hd__mux2_1 _15249_ (.A0(_02426_),
    .A1(\cur_mb_mem[68][0] ),
    .S(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__clkbuf_1 _15250_ (.A(_02463_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _15251_ (.A0(_02429_),
    .A1(net1600),
    .S(_02462_),
    .X(_02464_));
 sky130_fd_sc_hd__clkbuf_1 _15252_ (.A(_02464_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _15253_ (.A0(_02431_),
    .A1(\cur_mb_mem[68][2] ),
    .S(_02462_),
    .X(_02465_));
 sky130_fd_sc_hd__clkbuf_1 _15254_ (.A(_02465_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _15255_ (.A0(_02433_),
    .A1(\cur_mb_mem[68][3] ),
    .S(_02462_),
    .X(_02466_));
 sky130_fd_sc_hd__clkbuf_1 _15256_ (.A(_02466_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _15257_ (.A0(_02435_),
    .A1(net705),
    .S(_02462_),
    .X(_02467_));
 sky130_fd_sc_hd__clkbuf_1 _15258_ (.A(_02467_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _15259_ (.A0(_02437_),
    .A1(net879),
    .S(_02462_),
    .X(_02468_));
 sky130_fd_sc_hd__clkbuf_1 _15260_ (.A(_02468_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _15261_ (.A0(_02439_),
    .A1(\cur_mb_mem[68][6] ),
    .S(_02462_),
    .X(_02469_));
 sky130_fd_sc_hd__clkbuf_1 _15262_ (.A(_02469_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _15263_ (.A0(_02441_),
    .A1(\cur_mb_mem[68][7] ),
    .S(_02462_),
    .X(_02470_));
 sky130_fd_sc_hd__clkbuf_1 _15264_ (.A(_02470_),
    .X(_00702_));
 sky130_fd_sc_hd__nand2_8 _15265_ (.A(_06218_),
    .B(_02443_),
    .Y(_02471_));
 sky130_fd_sc_hd__mux2_1 _15266_ (.A0(_02426_),
    .A1(net723),
    .S(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__clkbuf_1 _15267_ (.A(_02472_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _15268_ (.A0(_02429_),
    .A1(net933),
    .S(_02471_),
    .X(_02473_));
 sky130_fd_sc_hd__clkbuf_1 _15269_ (.A(_02473_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _15270_ (.A0(_02431_),
    .A1(\cur_mb_mem[69][2] ),
    .S(_02471_),
    .X(_02474_));
 sky130_fd_sc_hd__clkbuf_1 _15271_ (.A(_02474_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _15272_ (.A0(_02433_),
    .A1(net1106),
    .S(_02471_),
    .X(_02475_));
 sky130_fd_sc_hd__clkbuf_1 _15273_ (.A(_02475_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _15274_ (.A0(_02435_),
    .A1(net1933),
    .S(_02471_),
    .X(_02476_));
 sky130_fd_sc_hd__clkbuf_1 _15275_ (.A(_02476_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _15276_ (.A0(_02437_),
    .A1(net1968),
    .S(_02471_),
    .X(_02477_));
 sky130_fd_sc_hd__clkbuf_1 _15277_ (.A(_02477_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _15278_ (.A0(_02439_),
    .A1(\cur_mb_mem[69][6] ),
    .S(_02471_),
    .X(_02478_));
 sky130_fd_sc_hd__clkbuf_1 _15279_ (.A(_02478_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _15280_ (.A0(_02441_),
    .A1(\cur_mb_mem[69][7] ),
    .S(_02471_),
    .X(_02479_));
 sky130_fd_sc_hd__clkbuf_1 _15281_ (.A(_02479_),
    .X(_00710_));
 sky130_fd_sc_hd__nand2_8 _15282_ (.A(_06144_),
    .B(_02443_),
    .Y(_02480_));
 sky130_fd_sc_hd__mux2_1 _15283_ (.A0(_02426_),
    .A1(net1091),
    .S(_02480_),
    .X(_02481_));
 sky130_fd_sc_hd__clkbuf_1 _15284_ (.A(_02481_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _15285_ (.A0(_02429_),
    .A1(\cur_mb_mem[70][1] ),
    .S(_02480_),
    .X(_02482_));
 sky130_fd_sc_hd__clkbuf_1 _15286_ (.A(_02482_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _15287_ (.A0(_02431_),
    .A1(net979),
    .S(_02480_),
    .X(_02483_));
 sky130_fd_sc_hd__clkbuf_1 _15288_ (.A(_02483_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _15289_ (.A0(_02433_),
    .A1(net1002),
    .S(_02480_),
    .X(_02484_));
 sky130_fd_sc_hd__clkbuf_1 _15290_ (.A(_02484_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _15291_ (.A0(_02435_),
    .A1(net1922),
    .S(_02480_),
    .X(_02485_));
 sky130_fd_sc_hd__clkbuf_1 _15292_ (.A(_02485_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _15293_ (.A0(_02437_),
    .A1(\cur_mb_mem[70][5] ),
    .S(_02480_),
    .X(_02486_));
 sky130_fd_sc_hd__clkbuf_1 _15294_ (.A(_02486_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _15295_ (.A0(_02439_),
    .A1(\cur_mb_mem[70][6] ),
    .S(_02480_),
    .X(_02487_));
 sky130_fd_sc_hd__clkbuf_1 _15296_ (.A(_02487_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _15297_ (.A0(_02441_),
    .A1(net1959),
    .S(_02480_),
    .X(_02488_));
 sky130_fd_sc_hd__clkbuf_1 _15298_ (.A(_02488_),
    .X(_00718_));
 sky130_fd_sc_hd__nand2_8 _15299_ (.A(_06460_),
    .B(_02443_),
    .Y(_02489_));
 sky130_fd_sc_hd__mux2_1 _15300_ (.A0(_02426_),
    .A1(net1529),
    .S(_02489_),
    .X(_02490_));
 sky130_fd_sc_hd__clkbuf_1 _15301_ (.A(_02490_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _15302_ (.A0(_02429_),
    .A1(\cur_mb_mem[71][1] ),
    .S(_02489_),
    .X(_02491_));
 sky130_fd_sc_hd__clkbuf_1 _15303_ (.A(_02491_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _15304_ (.A0(_02431_),
    .A1(net501),
    .S(_02489_),
    .X(_02492_));
 sky130_fd_sc_hd__clkbuf_1 _15305_ (.A(_02492_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _15306_ (.A0(_02433_),
    .A1(\cur_mb_mem[71][3] ),
    .S(_02489_),
    .X(_02493_));
 sky130_fd_sc_hd__clkbuf_1 _15307_ (.A(_02493_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _15308_ (.A0(_02435_),
    .A1(net737),
    .S(_02489_),
    .X(_02494_));
 sky130_fd_sc_hd__clkbuf_1 _15309_ (.A(_02494_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _15310_ (.A0(_02437_),
    .A1(net1281),
    .S(_02489_),
    .X(_02495_));
 sky130_fd_sc_hd__clkbuf_1 _15311_ (.A(_02495_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _15312_ (.A0(_02439_),
    .A1(\cur_mb_mem[71][6] ),
    .S(_02489_),
    .X(_02496_));
 sky130_fd_sc_hd__clkbuf_1 _15313_ (.A(_02496_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _15314_ (.A0(_02441_),
    .A1(\cur_mb_mem[71][7] ),
    .S(_02489_),
    .X(_02497_));
 sky130_fd_sc_hd__clkbuf_1 _15315_ (.A(_02497_),
    .X(_00726_));
 sky130_fd_sc_hd__nand2_8 _15316_ (.A(_06288_),
    .B(_02443_),
    .Y(_02498_));
 sky130_fd_sc_hd__mux2_1 _15317_ (.A0(_02426_),
    .A1(net1831),
    .S(_02498_),
    .X(_02499_));
 sky130_fd_sc_hd__clkbuf_1 _15318_ (.A(_02499_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _15319_ (.A0(_02429_),
    .A1(\cur_mb_mem[72][1] ),
    .S(_02498_),
    .X(_02500_));
 sky130_fd_sc_hd__clkbuf_1 _15320_ (.A(_02500_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _15321_ (.A0(_02431_),
    .A1(net1669),
    .S(_02498_),
    .X(_02501_));
 sky130_fd_sc_hd__clkbuf_1 _15322_ (.A(_02501_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _15323_ (.A0(_02433_),
    .A1(net404),
    .S(_02498_),
    .X(_02502_));
 sky130_fd_sc_hd__clkbuf_1 _15324_ (.A(_02502_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _15325_ (.A0(_02435_),
    .A1(net1228),
    .S(_02498_),
    .X(_02503_));
 sky130_fd_sc_hd__clkbuf_1 _15326_ (.A(_02503_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _15327_ (.A0(_02437_),
    .A1(net1332),
    .S(_02498_),
    .X(_02504_));
 sky130_fd_sc_hd__clkbuf_1 _15328_ (.A(_02504_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _15329_ (.A0(_02439_),
    .A1(net1368),
    .S(_02498_),
    .X(_02505_));
 sky130_fd_sc_hd__clkbuf_1 _15330_ (.A(_02505_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _15331_ (.A0(_02441_),
    .A1(net1030),
    .S(_02498_),
    .X(_02506_));
 sky130_fd_sc_hd__clkbuf_1 _15332_ (.A(_02506_),
    .X(_00734_));
 sky130_fd_sc_hd__nand2_8 _15333_ (.A(_06328_),
    .B(_02443_),
    .Y(_02507_));
 sky130_fd_sc_hd__mux2_1 _15334_ (.A0(_02426_),
    .A1(\cur_mb_mem[73][0] ),
    .S(_02507_),
    .X(_02508_));
 sky130_fd_sc_hd__clkbuf_1 _15335_ (.A(_02508_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _15336_ (.A0(_02429_),
    .A1(net909),
    .S(_02507_),
    .X(_02509_));
 sky130_fd_sc_hd__clkbuf_1 _15337_ (.A(_02509_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _15338_ (.A0(_02431_),
    .A1(net1986),
    .S(_02507_),
    .X(_02510_));
 sky130_fd_sc_hd__clkbuf_1 _15339_ (.A(_02510_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _15340_ (.A0(_02433_),
    .A1(\cur_mb_mem[73][3] ),
    .S(_02507_),
    .X(_02511_));
 sky130_fd_sc_hd__clkbuf_1 _15341_ (.A(_02511_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _15342_ (.A0(_02435_),
    .A1(\cur_mb_mem[73][4] ),
    .S(_02507_),
    .X(_02512_));
 sky130_fd_sc_hd__clkbuf_1 _15343_ (.A(_02512_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _15344_ (.A0(_02437_),
    .A1(\cur_mb_mem[73][5] ),
    .S(_02507_),
    .X(_02513_));
 sky130_fd_sc_hd__clkbuf_1 _15345_ (.A(_02513_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _15346_ (.A0(_02439_),
    .A1(\cur_mb_mem[73][6] ),
    .S(_02507_),
    .X(_02514_));
 sky130_fd_sc_hd__clkbuf_1 _15347_ (.A(_02514_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _15348_ (.A0(_02441_),
    .A1(\cur_mb_mem[73][7] ),
    .S(_02507_),
    .X(_02515_));
 sky130_fd_sc_hd__clkbuf_1 _15349_ (.A(_02515_),
    .X(_00742_));
 sky130_fd_sc_hd__nand2_8 _15350_ (.A(_06417_),
    .B(_02443_),
    .Y(_02516_));
 sky130_fd_sc_hd__mux2_1 _15351_ (.A0(_02426_),
    .A1(\cur_mb_mem[74][0] ),
    .S(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__clkbuf_1 _15352_ (.A(_02517_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _15353_ (.A0(_02429_),
    .A1(net1734),
    .S(_02516_),
    .X(_02518_));
 sky130_fd_sc_hd__clkbuf_1 _15354_ (.A(_02518_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _15355_ (.A0(_02431_),
    .A1(\cur_mb_mem[74][2] ),
    .S(_02516_),
    .X(_02519_));
 sky130_fd_sc_hd__clkbuf_1 _15356_ (.A(_02519_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _15357_ (.A0(_02433_),
    .A1(\cur_mb_mem[74][3] ),
    .S(_02516_),
    .X(_02520_));
 sky130_fd_sc_hd__clkbuf_1 _15358_ (.A(_02520_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _15359_ (.A0(_02435_),
    .A1(\cur_mb_mem[74][4] ),
    .S(_02516_),
    .X(_02521_));
 sky130_fd_sc_hd__clkbuf_1 _15360_ (.A(_02521_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _15361_ (.A0(_02437_),
    .A1(\cur_mb_mem[74][5] ),
    .S(_02516_),
    .X(_02522_));
 sky130_fd_sc_hd__clkbuf_1 _15362_ (.A(_02522_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _15363_ (.A0(_02439_),
    .A1(net1753),
    .S(_02516_),
    .X(_02523_));
 sky130_fd_sc_hd__clkbuf_1 _15364_ (.A(_02523_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _15365_ (.A0(_02441_),
    .A1(\cur_mb_mem[74][7] ),
    .S(_02516_),
    .X(_02524_));
 sky130_fd_sc_hd__clkbuf_1 _15366_ (.A(_02524_),
    .X(_00750_));
 sky130_fd_sc_hd__buf_6 _15367_ (.A(_09132_),
    .X(_02525_));
 sky130_fd_sc_hd__buf_8 _15368_ (.A(_06049_),
    .X(_02526_));
 sky130_fd_sc_hd__nand3_4 _15369_ (.A(_02526_),
    .B(_06024_),
    .C(_08901_),
    .Y(_02527_));
 sky130_fd_sc_hd__mux2_1 _15370_ (.A0(_02525_),
    .A1(net1362),
    .S(net218),
    .X(_02528_));
 sky130_fd_sc_hd__clkbuf_1 _15371_ (.A(_02528_),
    .X(_00751_));
 sky130_fd_sc_hd__buf_4 _15372_ (.A(_09136_),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _15373_ (.A0(_02529_),
    .A1(net1254),
    .S(_02527_),
    .X(_02530_));
 sky130_fd_sc_hd__clkbuf_1 _15374_ (.A(_02530_),
    .X(_00752_));
 sky130_fd_sc_hd__clkbuf_8 _15375_ (.A(_09139_),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _15376_ (.A0(_02531_),
    .A1(net939),
    .S(net218),
    .X(_02532_));
 sky130_fd_sc_hd__clkbuf_1 _15377_ (.A(_02532_),
    .X(_00753_));
 sky130_fd_sc_hd__clkbuf_8 _15378_ (.A(_09142_),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _15379_ (.A0(_02533_),
    .A1(net1526),
    .S(net218),
    .X(_02534_));
 sky130_fd_sc_hd__clkbuf_1 _15380_ (.A(_02534_),
    .X(_00754_));
 sky130_fd_sc_hd__buf_4 _15381_ (.A(_09145_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _15382_ (.A0(_02535_),
    .A1(net594),
    .S(_02527_),
    .X(_02536_));
 sky130_fd_sc_hd__clkbuf_1 _15383_ (.A(_02536_),
    .X(_00755_));
 sky130_fd_sc_hd__buf_4 _15384_ (.A(_09148_),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _15385_ (.A0(_02537_),
    .A1(net693),
    .S(_02527_),
    .X(_02538_));
 sky130_fd_sc_hd__clkbuf_1 _15386_ (.A(_02538_),
    .X(_00756_));
 sky130_fd_sc_hd__clkbuf_4 _15387_ (.A(_09151_),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _15388_ (.A0(_02539_),
    .A1(\cur_mb_mem[75][6] ),
    .S(_02527_),
    .X(_02540_));
 sky130_fd_sc_hd__clkbuf_1 _15389_ (.A(_02540_),
    .X(_00757_));
 sky130_fd_sc_hd__buf_4 _15390_ (.A(_09154_),
    .X(_02541_));
 sky130_fd_sc_hd__mux2_1 _15391_ (.A0(_02541_),
    .A1(net1107),
    .S(net218),
    .X(_02542_));
 sky130_fd_sc_hd__clkbuf_1 _15392_ (.A(_02542_),
    .X(_00758_));
 sky130_fd_sc_hd__nand2_8 _15393_ (.A(_06340_),
    .B(_02443_),
    .Y(_02543_));
 sky130_fd_sc_hd__mux2_1 _15394_ (.A0(_02525_),
    .A1(net617),
    .S(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__clkbuf_1 _15395_ (.A(_02544_),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _15396_ (.A0(_02529_),
    .A1(net1103),
    .S(_02543_),
    .X(_02545_));
 sky130_fd_sc_hd__clkbuf_1 _15397_ (.A(_02545_),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _15398_ (.A0(_02531_),
    .A1(net616),
    .S(_02543_),
    .X(_02546_));
 sky130_fd_sc_hd__clkbuf_1 _15399_ (.A(_02546_),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _15400_ (.A0(_02533_),
    .A1(net478),
    .S(_02543_),
    .X(_02547_));
 sky130_fd_sc_hd__clkbuf_1 _15401_ (.A(_02547_),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _15402_ (.A0(_02535_),
    .A1(net487),
    .S(_02543_),
    .X(_02548_));
 sky130_fd_sc_hd__clkbuf_1 _15403_ (.A(_02548_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _15404_ (.A0(_02537_),
    .A1(net685),
    .S(_02543_),
    .X(_02549_));
 sky130_fd_sc_hd__clkbuf_1 _15405_ (.A(_02549_),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _15406_ (.A0(_02539_),
    .A1(net1537),
    .S(_02543_),
    .X(_02550_));
 sky130_fd_sc_hd__clkbuf_1 _15407_ (.A(_02550_),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _15408_ (.A0(_02541_),
    .A1(\cur_mb_mem[76][7] ),
    .S(_02543_),
    .X(_02551_));
 sky130_fd_sc_hd__clkbuf_1 _15409_ (.A(_02551_),
    .X(_00766_));
 sky130_fd_sc_hd__buf_12 _15410_ (.A(_08958_),
    .X(_02552_));
 sky130_fd_sc_hd__nand2_8 _15411_ (.A(_06058_),
    .B(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__mux2_1 _15412_ (.A0(_02525_),
    .A1(net844),
    .S(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__clkbuf_1 _15413_ (.A(_02554_),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _15414_ (.A0(_02529_),
    .A1(net1532),
    .S(_02553_),
    .X(_02555_));
 sky130_fd_sc_hd__clkbuf_1 _15415_ (.A(_02555_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _15416_ (.A0(_02531_),
    .A1(net1909),
    .S(_02553_),
    .X(_02556_));
 sky130_fd_sc_hd__clkbuf_1 _15417_ (.A(_02556_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _15418_ (.A0(_02533_),
    .A1(net743),
    .S(_02553_),
    .X(_02557_));
 sky130_fd_sc_hd__clkbuf_1 _15419_ (.A(_02557_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _15420_ (.A0(_02535_),
    .A1(net655),
    .S(_02553_),
    .X(_02558_));
 sky130_fd_sc_hd__clkbuf_1 _15421_ (.A(_02558_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _15422_ (.A0(_02537_),
    .A1(net954),
    .S(_02553_),
    .X(_02559_));
 sky130_fd_sc_hd__clkbuf_1 _15423_ (.A(_02559_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _15424_ (.A0(_02539_),
    .A1(\cur_mb_mem[77][6] ),
    .S(_02553_),
    .X(_02560_));
 sky130_fd_sc_hd__clkbuf_1 _15425_ (.A(_02560_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _15426_ (.A0(_02541_),
    .A1(net1382),
    .S(_02553_),
    .X(_02561_));
 sky130_fd_sc_hd__clkbuf_1 _15427_ (.A(_02561_),
    .X(_00774_));
 sky130_fd_sc_hd__nand3_4 _15428_ (.A(_06024_),
    .B(_09036_),
    .C(_08901_),
    .Y(_02562_));
 sky130_fd_sc_hd__mux2_1 _15429_ (.A0(_02525_),
    .A1(net691),
    .S(_02562_),
    .X(_02563_));
 sky130_fd_sc_hd__clkbuf_1 _15430_ (.A(_02563_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _15431_ (.A0(_02529_),
    .A1(net1047),
    .S(_02562_),
    .X(_02564_));
 sky130_fd_sc_hd__clkbuf_1 _15432_ (.A(_02564_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _15433_ (.A0(_02531_),
    .A1(net1560),
    .S(_02562_),
    .X(_02565_));
 sky130_fd_sc_hd__clkbuf_1 _15434_ (.A(_02565_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _15435_ (.A0(_02533_),
    .A1(net847),
    .S(_02562_),
    .X(_02566_));
 sky130_fd_sc_hd__clkbuf_1 _15436_ (.A(_02566_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _15437_ (.A0(_02535_),
    .A1(net1004),
    .S(_02562_),
    .X(_02567_));
 sky130_fd_sc_hd__clkbuf_1 _15438_ (.A(_02567_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _15439_ (.A0(_02537_),
    .A1(net848),
    .S(_02562_),
    .X(_02568_));
 sky130_fd_sc_hd__clkbuf_1 _15440_ (.A(_02568_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _15441_ (.A0(_02539_),
    .A1(net861),
    .S(_02562_),
    .X(_02569_));
 sky130_fd_sc_hd__clkbuf_1 _15442_ (.A(_02569_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _15443_ (.A0(_02541_),
    .A1(net1413),
    .S(_02562_),
    .X(_02570_));
 sky130_fd_sc_hd__clkbuf_1 _15444_ (.A(_02570_),
    .X(_00782_));
 sky130_fd_sc_hd__nand2_8 _15445_ (.A(_06122_),
    .B(_02552_),
    .Y(_02571_));
 sky130_fd_sc_hd__mux2_1 _15446_ (.A0(_02525_),
    .A1(\cur_mb_mem[79][0] ),
    .S(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__clkbuf_1 _15447_ (.A(_02572_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _15448_ (.A0(_02529_),
    .A1(net961),
    .S(_02571_),
    .X(_02573_));
 sky130_fd_sc_hd__clkbuf_1 _15449_ (.A(_02573_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _15450_ (.A0(_02531_),
    .A1(\cur_mb_mem[79][2] ),
    .S(_02571_),
    .X(_02574_));
 sky130_fd_sc_hd__clkbuf_1 _15451_ (.A(_02574_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _15452_ (.A0(_02533_),
    .A1(\cur_mb_mem[79][3] ),
    .S(_02571_),
    .X(_02575_));
 sky130_fd_sc_hd__clkbuf_1 _15453_ (.A(_02575_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _15454_ (.A0(_02535_),
    .A1(net1890),
    .S(_02571_),
    .X(_02576_));
 sky130_fd_sc_hd__clkbuf_1 _15455_ (.A(_02576_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _15456_ (.A0(_02537_),
    .A1(\cur_mb_mem[79][5] ),
    .S(_02571_),
    .X(_02577_));
 sky130_fd_sc_hd__clkbuf_1 _15457_ (.A(_02577_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _15458_ (.A0(_02539_),
    .A1(net1347),
    .S(_02571_),
    .X(_02578_));
 sky130_fd_sc_hd__clkbuf_1 _15459_ (.A(_02578_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _15460_ (.A0(_02541_),
    .A1(\cur_mb_mem[79][7] ),
    .S(_02571_),
    .X(_02579_));
 sky130_fd_sc_hd__clkbuf_1 _15461_ (.A(_02579_),
    .X(_00790_));
 sky130_fd_sc_hd__buf_4 _15462_ (.A(_05916_),
    .X(_02580_));
 sky130_fd_sc_hd__nand2_8 _15463_ (.A(_02580_),
    .B(_08883_),
    .Y(_02581_));
 sky130_fd_sc_hd__mux2_1 _15464_ (.A0(_02525_),
    .A1(net531),
    .S(_02581_),
    .X(_02582_));
 sky130_fd_sc_hd__clkbuf_1 _15465_ (.A(_02582_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _15466_ (.A0(_02529_),
    .A1(\cur_mb_mem[80][1] ),
    .S(_02581_),
    .X(_02583_));
 sky130_fd_sc_hd__clkbuf_1 _15467_ (.A(_02583_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _15468_ (.A0(_02531_),
    .A1(net1169),
    .S(_02581_),
    .X(_02584_));
 sky130_fd_sc_hd__clkbuf_1 _15469_ (.A(_02584_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _15470_ (.A0(_02533_),
    .A1(net1130),
    .S(_02581_),
    .X(_02585_));
 sky130_fd_sc_hd__clkbuf_1 _15471_ (.A(_02585_),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _15472_ (.A0(_02535_),
    .A1(net1766),
    .S(_02581_),
    .X(_02586_));
 sky130_fd_sc_hd__clkbuf_1 _15473_ (.A(_02586_),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _15474_ (.A0(_02537_),
    .A1(net1711),
    .S(_02581_),
    .X(_02587_));
 sky130_fd_sc_hd__clkbuf_1 _15475_ (.A(_02587_),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _15476_ (.A0(_02539_),
    .A1(net1516),
    .S(_02581_),
    .X(_02588_));
 sky130_fd_sc_hd__clkbuf_1 _15477_ (.A(_02588_),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _15478_ (.A0(_02541_),
    .A1(\cur_mb_mem[80][7] ),
    .S(_02581_),
    .X(_02589_));
 sky130_fd_sc_hd__clkbuf_1 _15479_ (.A(_02589_),
    .X(_00798_));
 sky130_fd_sc_hd__or3_1 _15480_ (.A(_06296_),
    .B(_05963_),
    .C(_08532_),
    .X(_02590_));
 sky130_fd_sc_hd__buf_6 _15481_ (.A(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__mux2_1 _15482_ (.A0(_02525_),
    .A1(net653),
    .S(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__clkbuf_1 _15483_ (.A(_02592_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _15484_ (.A0(_02529_),
    .A1(net856),
    .S(_02591_),
    .X(_02593_));
 sky130_fd_sc_hd__clkbuf_1 _15485_ (.A(_02593_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _15486_ (.A0(_02531_),
    .A1(\cur_mb_mem[81][2] ),
    .S(_02591_),
    .X(_02594_));
 sky130_fd_sc_hd__clkbuf_1 _15487_ (.A(_02594_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _15488_ (.A0(_02533_),
    .A1(net1009),
    .S(_02591_),
    .X(_02595_));
 sky130_fd_sc_hd__clkbuf_1 _15489_ (.A(_02595_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _15490_ (.A0(_02535_),
    .A1(net1587),
    .S(_02591_),
    .X(_02596_));
 sky130_fd_sc_hd__clkbuf_1 _15491_ (.A(_02596_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _15492_ (.A0(_02537_),
    .A1(net905),
    .S(_02591_),
    .X(_02597_));
 sky130_fd_sc_hd__clkbuf_1 _15493_ (.A(_02597_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _15494_ (.A0(_02539_),
    .A1(net1317),
    .S(_02591_),
    .X(_02598_));
 sky130_fd_sc_hd__clkbuf_1 _15495_ (.A(_02598_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _15496_ (.A0(_02541_),
    .A1(\cur_mb_mem[81][7] ),
    .S(_02591_),
    .X(_02599_));
 sky130_fd_sc_hd__clkbuf_1 _15497_ (.A(_02599_),
    .X(_00806_));
 sky130_fd_sc_hd__or3_1 _15498_ (.A(_06265_),
    .B(_06296_),
    .C(_08532_),
    .X(_02600_));
 sky130_fd_sc_hd__clkbuf_8 _15499_ (.A(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__mux2_1 _15500_ (.A0(_02525_),
    .A1(net582),
    .S(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__clkbuf_1 _15501_ (.A(_02602_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _15502_ (.A0(_02529_),
    .A1(net872),
    .S(_02601_),
    .X(_02603_));
 sky130_fd_sc_hd__clkbuf_1 _15503_ (.A(_02603_),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _15504_ (.A0(_02531_),
    .A1(net679),
    .S(_02601_),
    .X(_02604_));
 sky130_fd_sc_hd__clkbuf_1 _15505_ (.A(_02604_),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_1 _15506_ (.A0(_02533_),
    .A1(net1054),
    .S(_02601_),
    .X(_02605_));
 sky130_fd_sc_hd__clkbuf_1 _15507_ (.A(_02605_),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _15508_ (.A0(_02535_),
    .A1(net924),
    .S(_02601_),
    .X(_02606_));
 sky130_fd_sc_hd__clkbuf_1 _15509_ (.A(_02606_),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _15510_ (.A0(_02537_),
    .A1(net613),
    .S(_02601_),
    .X(_02607_));
 sky130_fd_sc_hd__clkbuf_1 _15511_ (.A(_02607_),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_1 _15512_ (.A0(_02539_),
    .A1(net1206),
    .S(_02601_),
    .X(_02608_));
 sky130_fd_sc_hd__clkbuf_1 _15513_ (.A(_02608_),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _15514_ (.A0(_02541_),
    .A1(net987),
    .S(_02601_),
    .X(_02609_));
 sky130_fd_sc_hd__clkbuf_1 _15515_ (.A(_02609_),
    .X(_00814_));
 sky130_fd_sc_hd__and3_1 _15516_ (.A(_02580_),
    .B(_02266_),
    .C(_02395_),
    .X(_02610_));
 sky130_fd_sc_hd__buf_6 _15517_ (.A(_02610_),
    .X(_02611_));
 sky130_fd_sc_hd__mux2_1 _15518_ (.A0(net1746),
    .A1(_02328_),
    .S(_02611_),
    .X(_02612_));
 sky130_fd_sc_hd__clkbuf_1 _15519_ (.A(_02612_),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _15520_ (.A0(net1833),
    .A1(_02333_),
    .S(_02611_),
    .X(_02613_));
 sky130_fd_sc_hd__clkbuf_1 _15521_ (.A(_02613_),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _15522_ (.A0(net1580),
    .A1(_02336_),
    .S(_02611_),
    .X(_02614_));
 sky130_fd_sc_hd__clkbuf_1 _15523_ (.A(_02614_),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _15524_ (.A0(net1492),
    .A1(_02339_),
    .S(_02611_),
    .X(_02615_));
 sky130_fd_sc_hd__clkbuf_1 _15525_ (.A(_02615_),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _15526_ (.A0(net1870),
    .A1(_02342_),
    .S(_02611_),
    .X(_02616_));
 sky130_fd_sc_hd__clkbuf_1 _15527_ (.A(_02616_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _15528_ (.A0(net1748),
    .A1(_02345_),
    .S(_02611_),
    .X(_02617_));
 sky130_fd_sc_hd__clkbuf_1 _15529_ (.A(_02617_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _15530_ (.A0(net643),
    .A1(_02348_),
    .S(_02611_),
    .X(_02618_));
 sky130_fd_sc_hd__clkbuf_1 _15531_ (.A(_02618_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _15532_ (.A0(net567),
    .A1(_02351_),
    .S(_02611_),
    .X(_02619_));
 sky130_fd_sc_hd__clkbuf_1 _15533_ (.A(_02619_),
    .X(_00822_));
 sky130_fd_sc_hd__or3_1 _15534_ (.A(_06161_),
    .B(_06296_),
    .C(_08532_),
    .X(_02620_));
 sky130_fd_sc_hd__clkbuf_8 _15535_ (.A(_02620_),
    .X(_02621_));
 sky130_fd_sc_hd__mux2_1 _15536_ (.A0(_02525_),
    .A1(\cur_mb_mem[84][0] ),
    .S(_02621_),
    .X(_02622_));
 sky130_fd_sc_hd__clkbuf_1 _15537_ (.A(_02622_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _15538_ (.A0(_02529_),
    .A1(net778),
    .S(_02621_),
    .X(_02623_));
 sky130_fd_sc_hd__clkbuf_1 _15539_ (.A(_02623_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _15540_ (.A0(_02531_),
    .A1(net1865),
    .S(_02621_),
    .X(_02624_));
 sky130_fd_sc_hd__clkbuf_1 _15541_ (.A(_02624_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _15542_ (.A0(_02533_),
    .A1(net773),
    .S(_02621_),
    .X(_02625_));
 sky130_fd_sc_hd__clkbuf_1 _15543_ (.A(_02625_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _15544_ (.A0(_02535_),
    .A1(net708),
    .S(_02621_),
    .X(_02626_));
 sky130_fd_sc_hd__clkbuf_1 _15545_ (.A(_02626_),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _15546_ (.A0(_02537_),
    .A1(net802),
    .S(_02621_),
    .X(_02627_));
 sky130_fd_sc_hd__clkbuf_1 _15547_ (.A(_02627_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _15548_ (.A0(_02539_),
    .A1(\cur_mb_mem[84][6] ),
    .S(_02621_),
    .X(_02628_));
 sky130_fd_sc_hd__clkbuf_1 _15549_ (.A(_02628_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _15550_ (.A0(_02541_),
    .A1(net1288),
    .S(_02621_),
    .X(_02629_));
 sky130_fd_sc_hd__clkbuf_1 _15551_ (.A(_02629_),
    .X(_00830_));
 sky130_fd_sc_hd__and3_1 _15552_ (.A(_02580_),
    .B(_02286_),
    .C(_02395_),
    .X(_02630_));
 sky130_fd_sc_hd__clkbuf_8 _15553_ (.A(_02630_),
    .X(_02631_));
 sky130_fd_sc_hd__mux2_1 _15554_ (.A0(net1612),
    .A1(_02328_),
    .S(_02631_),
    .X(_02632_));
 sky130_fd_sc_hd__clkbuf_1 _15555_ (.A(_02632_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _15556_ (.A0(net807),
    .A1(_02333_),
    .S(_02631_),
    .X(_02633_));
 sky130_fd_sc_hd__clkbuf_1 _15557_ (.A(_02633_),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _15558_ (.A0(net1463),
    .A1(_02336_),
    .S(_02631_),
    .X(_02634_));
 sky130_fd_sc_hd__clkbuf_1 _15559_ (.A(_02634_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _15560_ (.A0(net762),
    .A1(_02339_),
    .S(_02631_),
    .X(_02635_));
 sky130_fd_sc_hd__clkbuf_1 _15561_ (.A(_02635_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _15562_ (.A0(net1512),
    .A1(_02342_),
    .S(_02631_),
    .X(_02636_));
 sky130_fd_sc_hd__clkbuf_1 _15563_ (.A(_02636_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _15564_ (.A0(net976),
    .A1(_02345_),
    .S(_02631_),
    .X(_02637_));
 sky130_fd_sc_hd__clkbuf_1 _15565_ (.A(_02637_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _15566_ (.A0(net1240),
    .A1(_02348_),
    .S(_02631_),
    .X(_02638_));
 sky130_fd_sc_hd__clkbuf_1 _15567_ (.A(_02638_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _15568_ (.A0(net588),
    .A1(_02351_),
    .S(_02631_),
    .X(_02639_));
 sky130_fd_sc_hd__clkbuf_1 _15569_ (.A(_02639_),
    .X(_00838_));
 sky130_fd_sc_hd__and3_1 _15570_ (.A(_02580_),
    .B(_02297_),
    .C(_02395_),
    .X(_02640_));
 sky130_fd_sc_hd__buf_6 _15571_ (.A(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__mux2_1 _15572_ (.A0(net364),
    .A1(_02328_),
    .S(_02641_),
    .X(_02642_));
 sky130_fd_sc_hd__clkbuf_1 _15573_ (.A(_02642_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _15574_ (.A0(net459),
    .A1(_02333_),
    .S(_02641_),
    .X(_02643_));
 sky130_fd_sc_hd__clkbuf_1 _15575_ (.A(_02643_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _15576_ (.A0(net1249),
    .A1(_02336_),
    .S(_02641_),
    .X(_02644_));
 sky130_fd_sc_hd__clkbuf_1 _15577_ (.A(_02644_),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _15578_ (.A0(net315),
    .A1(_02339_),
    .S(_02641_),
    .X(_02645_));
 sky130_fd_sc_hd__clkbuf_1 _15579_ (.A(_02645_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _15580_ (.A0(net572),
    .A1(_02342_),
    .S(_02641_),
    .X(_02646_));
 sky130_fd_sc_hd__clkbuf_1 _15581_ (.A(_02646_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _15582_ (.A0(net322),
    .A1(_02345_),
    .S(_02641_),
    .X(_02647_));
 sky130_fd_sc_hd__clkbuf_1 _15583_ (.A(_02647_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _15584_ (.A0(net884),
    .A1(_02348_),
    .S(_02641_),
    .X(_02648_));
 sky130_fd_sc_hd__clkbuf_1 _15585_ (.A(_02648_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _15586_ (.A0(net1077),
    .A1(_02351_),
    .S(_02641_),
    .X(_02649_));
 sky130_fd_sc_hd__clkbuf_1 _15587_ (.A(_02649_),
    .X(_00846_));
 sky130_fd_sc_hd__buf_12 _15588_ (.A(_02327_),
    .X(_02650_));
 sky130_fd_sc_hd__and3_1 _15589_ (.A(_02580_),
    .B(_08839_),
    .C(_02395_),
    .X(_02651_));
 sky130_fd_sc_hd__buf_8 _15590_ (.A(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__mux2_1 _15591_ (.A0(net578),
    .A1(_02650_),
    .S(_02652_),
    .X(_02653_));
 sky130_fd_sc_hd__clkbuf_1 _15592_ (.A(_02653_),
    .X(_00847_));
 sky130_fd_sc_hd__buf_6 _15593_ (.A(_02332_),
    .X(_02654_));
 sky130_fd_sc_hd__mux2_1 _15594_ (.A0(net373),
    .A1(_02654_),
    .S(_02652_),
    .X(_02655_));
 sky130_fd_sc_hd__clkbuf_1 _15595_ (.A(_02655_),
    .X(_00848_));
 sky130_fd_sc_hd__buf_12 _15596_ (.A(_02335_),
    .X(_02656_));
 sky130_fd_sc_hd__mux2_1 _15597_ (.A0(net425),
    .A1(_02656_),
    .S(_02652_),
    .X(_02657_));
 sky130_fd_sc_hd__clkbuf_1 _15598_ (.A(_02657_),
    .X(_00849_));
 sky130_fd_sc_hd__buf_12 _15599_ (.A(_02338_),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _15600_ (.A0(net347),
    .A1(_02658_),
    .S(_02652_),
    .X(_02659_));
 sky130_fd_sc_hd__clkbuf_1 _15601_ (.A(_02659_),
    .X(_00850_));
 sky130_fd_sc_hd__buf_6 _15602_ (.A(_02341_),
    .X(_02660_));
 sky130_fd_sc_hd__mux2_1 _15603_ (.A0(net360),
    .A1(_02660_),
    .S(_02652_),
    .X(_02661_));
 sky130_fd_sc_hd__clkbuf_1 _15604_ (.A(_02661_),
    .X(_00851_));
 sky130_fd_sc_hd__buf_6 _15605_ (.A(_02344_),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _15606_ (.A0(net554),
    .A1(_02662_),
    .S(_02652_),
    .X(_02663_));
 sky130_fd_sc_hd__clkbuf_1 _15607_ (.A(_02663_),
    .X(_00852_));
 sky130_fd_sc_hd__buf_4 _15608_ (.A(_02347_),
    .X(_02664_));
 sky130_fd_sc_hd__mux2_1 _15609_ (.A0(net850),
    .A1(_02664_),
    .S(_02652_),
    .X(_02665_));
 sky130_fd_sc_hd__clkbuf_1 _15610_ (.A(_02665_),
    .X(_00853_));
 sky130_fd_sc_hd__buf_4 _15611_ (.A(_02350_),
    .X(_02666_));
 sky130_fd_sc_hd__mux2_1 _15612_ (.A0(net1506),
    .A1(_02666_),
    .S(_02652_),
    .X(_02667_));
 sky130_fd_sc_hd__clkbuf_1 _15613_ (.A(_02667_),
    .X(_00854_));
 sky130_fd_sc_hd__or3_1 _15614_ (.A(_06276_),
    .B(_06296_),
    .C(_08532_),
    .X(_02668_));
 sky130_fd_sc_hd__buf_4 _15615_ (.A(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__mux2_1 _15616_ (.A0(_02525_),
    .A1(net1892),
    .S(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__clkbuf_1 _15617_ (.A(_02670_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _15618_ (.A0(_02529_),
    .A1(\cur_mb_mem[88][1] ),
    .S(_02669_),
    .X(_02671_));
 sky130_fd_sc_hd__clkbuf_1 _15619_ (.A(_02671_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _15620_ (.A0(_02531_),
    .A1(net985),
    .S(_02669_),
    .X(_02672_));
 sky130_fd_sc_hd__clkbuf_1 _15621_ (.A(_02672_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _15622_ (.A0(_02533_),
    .A1(net877),
    .S(_02669_),
    .X(_02673_));
 sky130_fd_sc_hd__clkbuf_1 _15623_ (.A(_02673_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _15624_ (.A0(_02535_),
    .A1(net741),
    .S(_02669_),
    .X(_02674_));
 sky130_fd_sc_hd__clkbuf_1 _15625_ (.A(_02674_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _15626_ (.A0(_02537_),
    .A1(net645),
    .S(_02669_),
    .X(_02675_));
 sky130_fd_sc_hd__clkbuf_1 _15627_ (.A(_02675_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _15628_ (.A0(_02539_),
    .A1(net1617),
    .S(_02669_),
    .X(_02676_));
 sky130_fd_sc_hd__clkbuf_1 _15629_ (.A(_02676_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _15630_ (.A0(_02541_),
    .A1(net1358),
    .S(_02669_),
    .X(_02677_));
 sky130_fd_sc_hd__clkbuf_1 _15631_ (.A(_02677_),
    .X(_00862_));
 sky130_fd_sc_hd__and3_1 _15632_ (.A(_08978_),
    .B(_02580_),
    .C(_02395_),
    .X(_02678_));
 sky130_fd_sc_hd__buf_4 _15633_ (.A(_02678_),
    .X(_02679_));
 sky130_fd_sc_hd__mux2_1 _15634_ (.A0(net346),
    .A1(_02650_),
    .S(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__clkbuf_1 _15635_ (.A(_02680_),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _15636_ (.A0(net336),
    .A1(_02654_),
    .S(_02679_),
    .X(_02681_));
 sky130_fd_sc_hd__clkbuf_1 _15637_ (.A(_02681_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _15638_ (.A0(net917),
    .A1(_02656_),
    .S(_02679_),
    .X(_02682_));
 sky130_fd_sc_hd__clkbuf_1 _15639_ (.A(_02682_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _15640_ (.A0(net311),
    .A1(_02658_),
    .S(_02679_),
    .X(_02683_));
 sky130_fd_sc_hd__clkbuf_1 _15641_ (.A(_02683_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _15642_ (.A0(net465),
    .A1(_02660_),
    .S(_02679_),
    .X(_02684_));
 sky130_fd_sc_hd__clkbuf_1 _15643_ (.A(_02684_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _15644_ (.A0(net517),
    .A1(_02662_),
    .S(_02679_),
    .X(_02685_));
 sky130_fd_sc_hd__clkbuf_1 _15645_ (.A(_02685_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _15646_ (.A0(net1328),
    .A1(_02664_),
    .S(_02679_),
    .X(_02686_));
 sky130_fd_sc_hd__clkbuf_1 _15647_ (.A(_02686_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _15648_ (.A0(net937),
    .A1(_02666_),
    .S(_02679_),
    .X(_02687_));
 sky130_fd_sc_hd__clkbuf_1 _15649_ (.A(_02687_),
    .X(_00870_));
 sky130_fd_sc_hd__and3_1 _15650_ (.A(_02353_),
    .B(_02580_),
    .C(_02395_),
    .X(_02688_));
 sky130_fd_sc_hd__buf_8 _15651_ (.A(_02688_),
    .X(_02689_));
 sky130_fd_sc_hd__mux2_1 _15652_ (.A0(net369),
    .A1(_02650_),
    .S(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__clkbuf_1 _15653_ (.A(_02690_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _15654_ (.A0(net823),
    .A1(_02654_),
    .S(_02689_),
    .X(_02691_));
 sky130_fd_sc_hd__clkbuf_1 _15655_ (.A(_02691_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _15656_ (.A0(net493),
    .A1(_02656_),
    .S(_02689_),
    .X(_02692_));
 sky130_fd_sc_hd__clkbuf_1 _15657_ (.A(_02692_),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _15658_ (.A0(net454),
    .A1(_02658_),
    .S(_02689_),
    .X(_02693_));
 sky130_fd_sc_hd__clkbuf_1 _15659_ (.A(_02693_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _15660_ (.A0(net755),
    .A1(_02660_),
    .S(_02689_),
    .X(_02694_));
 sky130_fd_sc_hd__clkbuf_1 _15661_ (.A(_02694_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _15662_ (.A0(net376),
    .A1(_02662_),
    .S(_02689_),
    .X(_02695_));
 sky130_fd_sc_hd__clkbuf_1 _15663_ (.A(_02695_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _15664_ (.A0(net1339),
    .A1(_02664_),
    .S(_02689_),
    .X(_02696_));
 sky130_fd_sc_hd__clkbuf_1 _15665_ (.A(_02696_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _15666_ (.A0(net381),
    .A1(_02666_),
    .S(_02689_),
    .X(_02697_));
 sky130_fd_sc_hd__clkbuf_1 _15667_ (.A(_02697_),
    .X(_00878_));
 sky130_fd_sc_hd__and3_1 _15668_ (.A(_02526_),
    .B(_02580_),
    .C(_02395_),
    .X(_02698_));
 sky130_fd_sc_hd__buf_8 _15669_ (.A(_02698_),
    .X(_02699_));
 sky130_fd_sc_hd__mux2_1 _15670_ (.A0(net871),
    .A1(_02650_),
    .S(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__clkbuf_1 _15671_ (.A(_02700_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _15672_ (.A0(net1607),
    .A1(_02654_),
    .S(_02699_),
    .X(_02701_));
 sky130_fd_sc_hd__clkbuf_1 _15673_ (.A(_02701_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _15674_ (.A0(net934),
    .A1(_02656_),
    .S(_02699_),
    .X(_02702_));
 sky130_fd_sc_hd__clkbuf_1 _15675_ (.A(_02702_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _15676_ (.A0(net766),
    .A1(_02658_),
    .S(_02699_),
    .X(_02703_));
 sky130_fd_sc_hd__clkbuf_1 _15677_ (.A(_02703_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _15678_ (.A0(net557),
    .A1(_02660_),
    .S(_02699_),
    .X(_02704_));
 sky130_fd_sc_hd__clkbuf_1 _15679_ (.A(_02704_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _15680_ (.A0(net488),
    .A1(_02662_),
    .S(_02699_),
    .X(_02705_));
 sky130_fd_sc_hd__clkbuf_1 _15681_ (.A(_02705_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _15682_ (.A0(net796),
    .A1(_02664_),
    .S(_02699_),
    .X(_02706_));
 sky130_fd_sc_hd__clkbuf_1 _15683_ (.A(_02706_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _15684_ (.A0(net622),
    .A1(_02666_),
    .S(_02699_),
    .X(_02707_));
 sky130_fd_sc_hd__clkbuf_1 _15685_ (.A(_02707_),
    .X(_00886_));
 sky130_fd_sc_hd__and3_1 _15686_ (.A(_02374_),
    .B(_05916_),
    .C(_02395_),
    .X(_02708_));
 sky130_fd_sc_hd__buf_8 _15687_ (.A(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__mux2_1 _15688_ (.A0(net491),
    .A1(_02650_),
    .S(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__clkbuf_1 _15689_ (.A(_02710_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _15690_ (.A0(net585),
    .A1(_02654_),
    .S(_02709_),
    .X(_02711_));
 sky130_fd_sc_hd__clkbuf_1 _15691_ (.A(_02711_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _15692_ (.A0(net494),
    .A1(_02656_),
    .S(_02709_),
    .X(_02712_));
 sky130_fd_sc_hd__clkbuf_1 _15693_ (.A(_02712_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _15694_ (.A0(net497),
    .A1(_02658_),
    .S(_02709_),
    .X(_02713_));
 sky130_fd_sc_hd__clkbuf_1 _15695_ (.A(_02713_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _15696_ (.A0(net489),
    .A1(_02660_),
    .S(_02709_),
    .X(_02714_));
 sky130_fd_sc_hd__clkbuf_1 _15697_ (.A(_02714_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _15698_ (.A0(net466),
    .A1(_02662_),
    .S(_02709_),
    .X(_02715_));
 sky130_fd_sc_hd__clkbuf_1 _15699_ (.A(_02715_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _15700_ (.A0(net378),
    .A1(_02664_),
    .S(_02709_),
    .X(_02716_));
 sky130_fd_sc_hd__clkbuf_1 _15701_ (.A(_02716_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _15702_ (.A0(net356),
    .A1(_02666_),
    .S(_02709_),
    .X(_02717_));
 sky130_fd_sc_hd__clkbuf_1 _15703_ (.A(_02717_),
    .X(_00894_));
 sky130_fd_sc_hd__buf_2 _15704_ (.A(_08900_),
    .X(_02718_));
 sky130_fd_sc_hd__and3_1 _15705_ (.A(_02580_),
    .B(_09025_),
    .C(_02718_),
    .X(_02719_));
 sky130_fd_sc_hd__buf_8 _15706_ (.A(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__mux2_1 _15707_ (.A0(net317),
    .A1(_02650_),
    .S(_02720_),
    .X(_02721_));
 sky130_fd_sc_hd__clkbuf_1 _15708_ (.A(_02721_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _15709_ (.A0(net434),
    .A1(_02654_),
    .S(_02720_),
    .X(_02722_));
 sky130_fd_sc_hd__clkbuf_1 _15710_ (.A(_02722_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _15711_ (.A0(net392),
    .A1(_02656_),
    .S(_02720_),
    .X(_02723_));
 sky130_fd_sc_hd__clkbuf_1 _15712_ (.A(_02723_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _15713_ (.A0(net354),
    .A1(_02658_),
    .S(_02720_),
    .X(_02724_));
 sky130_fd_sc_hd__clkbuf_1 _15714_ (.A(_02724_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _15715_ (.A0(net332),
    .A1(_02660_),
    .S(_02720_),
    .X(_02725_));
 sky130_fd_sc_hd__clkbuf_1 _15716_ (.A(_02725_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _15717_ (.A0(net475),
    .A1(_02662_),
    .S(_02720_),
    .X(_02726_));
 sky130_fd_sc_hd__clkbuf_1 _15718_ (.A(_02726_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _15719_ (.A0(net362),
    .A1(_02664_),
    .S(_02720_),
    .X(_02727_));
 sky130_fd_sc_hd__clkbuf_1 _15720_ (.A(_02727_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _15721_ (.A0(net1066),
    .A1(_02666_),
    .S(_02720_),
    .X(_02728_));
 sky130_fd_sc_hd__clkbuf_1 _15722_ (.A(_02728_),
    .X(_00902_));
 sky130_fd_sc_hd__and3_1 _15723_ (.A(_02580_),
    .B(_09036_),
    .C(_02718_),
    .X(_02729_));
 sky130_fd_sc_hd__buf_8 _15724_ (.A(_02729_),
    .X(_02730_));
 sky130_fd_sc_hd__mux2_1 _15725_ (.A0(net507),
    .A1(_02650_),
    .S(_02730_),
    .X(_02731_));
 sky130_fd_sc_hd__clkbuf_1 _15726_ (.A(_02731_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _15727_ (.A0(net541),
    .A1(_02654_),
    .S(_02730_),
    .X(_02732_));
 sky130_fd_sc_hd__clkbuf_1 _15728_ (.A(_02732_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _15729_ (.A0(net553),
    .A1(_02656_),
    .S(_02730_),
    .X(_02733_));
 sky130_fd_sc_hd__clkbuf_1 _15730_ (.A(_02733_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _15731_ (.A0(net427),
    .A1(_02658_),
    .S(_02730_),
    .X(_02734_));
 sky130_fd_sc_hd__clkbuf_1 _15732_ (.A(_02734_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _15733_ (.A0(net558),
    .A1(_02660_),
    .S(_02730_),
    .X(_02735_));
 sky130_fd_sc_hd__clkbuf_1 _15734_ (.A(_02735_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _15735_ (.A0(net631),
    .A1(_02662_),
    .S(_02730_),
    .X(_02736_));
 sky130_fd_sc_hd__clkbuf_1 _15736_ (.A(_02736_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _15737_ (.A0(net735),
    .A1(_02664_),
    .S(_02730_),
    .X(_02737_));
 sky130_fd_sc_hd__clkbuf_1 _15738_ (.A(_02737_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _15739_ (.A0(net1023),
    .A1(_02666_),
    .S(_02730_),
    .X(_02738_));
 sky130_fd_sc_hd__clkbuf_1 _15740_ (.A(_02738_),
    .X(_00910_));
 sky130_fd_sc_hd__and3_1 _15741_ (.A(_02406_),
    .B(_05916_),
    .C(_02718_),
    .X(_02739_));
 sky130_fd_sc_hd__clkbuf_8 _15742_ (.A(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__mux2_1 _15743_ (.A0(net1141),
    .A1(_02650_),
    .S(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__clkbuf_1 _15744_ (.A(_02741_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _15745_ (.A0(net1340),
    .A1(_02654_),
    .S(_02740_),
    .X(_02742_));
 sky130_fd_sc_hd__clkbuf_1 _15746_ (.A(_02742_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _15747_ (.A0(net900),
    .A1(_02656_),
    .S(_02740_),
    .X(_02743_));
 sky130_fd_sc_hd__clkbuf_1 _15748_ (.A(_02743_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _15749_ (.A0(net1407),
    .A1(_02658_),
    .S(_02740_),
    .X(_02744_));
 sky130_fd_sc_hd__clkbuf_1 _15750_ (.A(_02744_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _15751_ (.A0(net490),
    .A1(_02660_),
    .S(_02740_),
    .X(_02745_));
 sky130_fd_sc_hd__clkbuf_1 _15752_ (.A(_02745_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _15753_ (.A0(net809),
    .A1(_02662_),
    .S(_02740_),
    .X(_02746_));
 sky130_fd_sc_hd__clkbuf_1 _15754_ (.A(_02746_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _15755_ (.A0(net883),
    .A1(_02664_),
    .S(_02740_),
    .X(_02747_));
 sky130_fd_sc_hd__clkbuf_1 _15756_ (.A(_02747_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _15757_ (.A0(net1383),
    .A1(_02666_),
    .S(_02740_),
    .X(_02748_));
 sky130_fd_sc_hd__clkbuf_1 _15758_ (.A(_02748_),
    .X(_00918_));
 sky130_fd_sc_hd__clkbuf_4 _15759_ (.A(_09132_),
    .X(_02749_));
 sky130_fd_sc_hd__buf_2 _15760_ (.A(_06299_),
    .X(_02750_));
 sky130_fd_sc_hd__nand2_4 _15761_ (.A(_02750_),
    .B(_08883_),
    .Y(_02751_));
 sky130_fd_sc_hd__mux2_1 _15762_ (.A0(_02749_),
    .A1(net1953),
    .S(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__clkbuf_1 _15763_ (.A(_02752_),
    .X(_00919_));
 sky130_fd_sc_hd__clkbuf_4 _15764_ (.A(_09136_),
    .X(_02753_));
 sky130_fd_sc_hd__mux2_1 _15765_ (.A0(_02753_),
    .A1(net1557),
    .S(_02751_),
    .X(_02754_));
 sky130_fd_sc_hd__clkbuf_1 _15766_ (.A(_02754_),
    .X(_00920_));
 sky130_fd_sc_hd__clkbuf_4 _15767_ (.A(_09139_),
    .X(_02755_));
 sky130_fd_sc_hd__mux2_1 _15768_ (.A0(_02755_),
    .A1(net1913),
    .S(_02751_),
    .X(_02756_));
 sky130_fd_sc_hd__clkbuf_1 _15769_ (.A(_02756_),
    .X(_00921_));
 sky130_fd_sc_hd__clkbuf_4 _15770_ (.A(_09142_),
    .X(_02757_));
 sky130_fd_sc_hd__mux2_1 _15771_ (.A0(_02757_),
    .A1(\cur_mb_mem[96][3] ),
    .S(_02751_),
    .X(_02758_));
 sky130_fd_sc_hd__clkbuf_1 _15772_ (.A(_02758_),
    .X(_00922_));
 sky130_fd_sc_hd__buf_4 _15773_ (.A(_09145_),
    .X(_02759_));
 sky130_fd_sc_hd__mux2_1 _15774_ (.A0(_02759_),
    .A1(net1954),
    .S(_02751_),
    .X(_02760_));
 sky130_fd_sc_hd__clkbuf_1 _15775_ (.A(_02760_),
    .X(_00923_));
 sky130_fd_sc_hd__clkbuf_4 _15776_ (.A(_09148_),
    .X(_02761_));
 sky130_fd_sc_hd__mux2_1 _15777_ (.A0(_02761_),
    .A1(net1911),
    .S(_02751_),
    .X(_02762_));
 sky130_fd_sc_hd__clkbuf_1 _15778_ (.A(_02762_),
    .X(_00924_));
 sky130_fd_sc_hd__clkbuf_4 _15779_ (.A(_09151_),
    .X(_02763_));
 sky130_fd_sc_hd__mux2_1 _15780_ (.A0(_02763_),
    .A1(\cur_mb_mem[96][6] ),
    .S(_02751_),
    .X(_02764_));
 sky130_fd_sc_hd__clkbuf_1 _15781_ (.A(_02764_),
    .X(_00925_));
 sky130_fd_sc_hd__clkbuf_4 _15782_ (.A(_09154_),
    .X(_02765_));
 sky130_fd_sc_hd__mux2_1 _15783_ (.A0(_02765_),
    .A1(\cur_mb_mem[96][7] ),
    .S(_02751_),
    .X(_02766_));
 sky130_fd_sc_hd__clkbuf_1 _15784_ (.A(_02766_),
    .X(_00926_));
 sky130_fd_sc_hd__nand2_4 _15785_ (.A(_06077_),
    .B(_02552_),
    .Y(_02767_));
 sky130_fd_sc_hd__mux2_1 _15786_ (.A0(_02749_),
    .A1(net1789),
    .S(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__clkbuf_1 _15787_ (.A(_02768_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _15788_ (.A0(_02753_),
    .A1(\cur_mb_mem[97][1] ),
    .S(_02767_),
    .X(_02769_));
 sky130_fd_sc_hd__clkbuf_1 _15789_ (.A(_02769_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _15790_ (.A0(_02755_),
    .A1(net1949),
    .S(_02767_),
    .X(_02770_));
 sky130_fd_sc_hd__clkbuf_1 _15791_ (.A(_02770_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _15792_ (.A0(_02757_),
    .A1(net1719),
    .S(_02767_),
    .X(_02771_));
 sky130_fd_sc_hd__clkbuf_1 _15793_ (.A(_02771_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _15794_ (.A0(_02759_),
    .A1(\cur_mb_mem[97][4] ),
    .S(_02767_),
    .X(_02772_));
 sky130_fd_sc_hd__clkbuf_1 _15795_ (.A(_02772_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _15796_ (.A0(_02761_),
    .A1(\cur_mb_mem[97][5] ),
    .S(_02767_),
    .X(_02773_));
 sky130_fd_sc_hd__clkbuf_1 _15797_ (.A(_02773_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _15798_ (.A0(_02763_),
    .A1(net1800),
    .S(_02767_),
    .X(_02774_));
 sky130_fd_sc_hd__clkbuf_1 _15799_ (.A(_02774_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _15800_ (.A0(_02765_),
    .A1(\cur_mb_mem[97][7] ),
    .S(_02767_),
    .X(_02775_));
 sky130_fd_sc_hd__clkbuf_1 _15801_ (.A(_02775_),
    .X(_00934_));
 sky130_fd_sc_hd__nand2_8 _15802_ (.A(_06330_),
    .B(_02552_),
    .Y(_02776_));
 sky130_fd_sc_hd__mux2_1 _15803_ (.A0(_02749_),
    .A1(\cur_mb_mem[98][0] ),
    .S(_02776_),
    .X(_02777_));
 sky130_fd_sc_hd__clkbuf_1 _15804_ (.A(_02777_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _15805_ (.A0(_02753_),
    .A1(\cur_mb_mem[98][1] ),
    .S(_02776_),
    .X(_02778_));
 sky130_fd_sc_hd__clkbuf_1 _15806_ (.A(_02778_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _15807_ (.A0(_02755_),
    .A1(\cur_mb_mem[98][2] ),
    .S(_02776_),
    .X(_02779_));
 sky130_fd_sc_hd__clkbuf_1 _15808_ (.A(_02779_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _15809_ (.A0(_02757_),
    .A1(\cur_mb_mem[98][3] ),
    .S(_02776_),
    .X(_02780_));
 sky130_fd_sc_hd__clkbuf_1 _15810_ (.A(_02780_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _15811_ (.A0(_02759_),
    .A1(\cur_mb_mem[98][4] ),
    .S(_02776_),
    .X(_02781_));
 sky130_fd_sc_hd__clkbuf_1 _15812_ (.A(_02781_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _15813_ (.A0(_02761_),
    .A1(\cur_mb_mem[98][5] ),
    .S(_02776_),
    .X(_02782_));
 sky130_fd_sc_hd__clkbuf_1 _15814_ (.A(_02782_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _15815_ (.A0(_02763_),
    .A1(\cur_mb_mem[98][6] ),
    .S(_02776_),
    .X(_02783_));
 sky130_fd_sc_hd__clkbuf_1 _15816_ (.A(_02783_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _15817_ (.A0(_02765_),
    .A1(\cur_mb_mem[98][7] ),
    .S(_02776_),
    .X(_02784_));
 sky130_fd_sc_hd__clkbuf_1 _15818_ (.A(_02784_),
    .X(_00942_));
 sky130_fd_sc_hd__and3_1 _15819_ (.A(_02750_),
    .B(_02266_),
    .C(_02718_),
    .X(_02785_));
 sky130_fd_sc_hd__buf_6 _15820_ (.A(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _15821_ (.A0(net527),
    .A1(_02650_),
    .S(_02786_),
    .X(_02787_));
 sky130_fd_sc_hd__clkbuf_1 _15822_ (.A(_02787_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _15823_ (.A0(net587),
    .A1(_02654_),
    .S(_02786_),
    .X(_02788_));
 sky130_fd_sc_hd__clkbuf_1 _15824_ (.A(_02788_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _15825_ (.A0(net528),
    .A1(_02656_),
    .S(_02786_),
    .X(_02789_));
 sky130_fd_sc_hd__clkbuf_1 _15826_ (.A(_02789_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _15827_ (.A0(net452),
    .A1(_02658_),
    .S(_02786_),
    .X(_02790_));
 sky130_fd_sc_hd__clkbuf_1 _15828_ (.A(_02790_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _15829_ (.A0(net457),
    .A1(_02660_),
    .S(_02786_),
    .X(_02791_));
 sky130_fd_sc_hd__clkbuf_1 _15830_ (.A(_02791_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _15831_ (.A0(net374),
    .A1(_02662_),
    .S(_02786_),
    .X(_02792_));
 sky130_fd_sc_hd__clkbuf_1 _15832_ (.A(_02792_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _15833_ (.A0(net891),
    .A1(_02664_),
    .S(_02786_),
    .X(_02793_));
 sky130_fd_sc_hd__clkbuf_1 _15834_ (.A(_02793_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _15835_ (.A0(net910),
    .A1(_02666_),
    .S(_02786_),
    .X(_02794_));
 sky130_fd_sc_hd__clkbuf_1 _15836_ (.A(_02794_),
    .X(_00950_));
 sky130_fd_sc_hd__nand2_4 _15837_ (.A(_06028_),
    .B(_02552_),
    .Y(_02795_));
 sky130_fd_sc_hd__mux2_1 _15838_ (.A0(_02749_),
    .A1(\cur_mb_mem[100][0] ),
    .S(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__clkbuf_1 _15839_ (.A(_02796_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _15840_ (.A0(_02753_),
    .A1(\cur_mb_mem[100][1] ),
    .S(_02795_),
    .X(_02797_));
 sky130_fd_sc_hd__clkbuf_1 _15841_ (.A(_02797_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _15842_ (.A0(_02755_),
    .A1(\cur_mb_mem[100][2] ),
    .S(_02795_),
    .X(_02798_));
 sky130_fd_sc_hd__clkbuf_1 _15843_ (.A(_02798_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _15844_ (.A0(_02757_),
    .A1(\cur_mb_mem[100][3] ),
    .S(_02795_),
    .X(_02799_));
 sky130_fd_sc_hd__clkbuf_1 _15845_ (.A(_02799_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _15846_ (.A0(_02759_),
    .A1(net1979),
    .S(_02795_),
    .X(_02800_));
 sky130_fd_sc_hd__clkbuf_1 _15847_ (.A(_02800_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _15848_ (.A0(_02761_),
    .A1(net1884),
    .S(_02795_),
    .X(_02801_));
 sky130_fd_sc_hd__clkbuf_1 _15849_ (.A(_02801_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _15850_ (.A0(_02763_),
    .A1(\cur_mb_mem[100][6] ),
    .S(_02795_),
    .X(_02802_));
 sky130_fd_sc_hd__clkbuf_1 _15851_ (.A(_02802_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _15852_ (.A0(_02765_),
    .A1(\cur_mb_mem[100][7] ),
    .S(_02795_),
    .X(_02803_));
 sky130_fd_sc_hd__clkbuf_1 _15853_ (.A(_02803_),
    .X(_00958_));
 sky130_fd_sc_hd__and3_1 _15854_ (.A(_02750_),
    .B(_02286_),
    .C(_02718_),
    .X(_02804_));
 sky130_fd_sc_hd__buf_8 _15855_ (.A(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_1 _15856_ (.A0(net886),
    .A1(_02650_),
    .S(_02805_),
    .X(_02806_));
 sky130_fd_sc_hd__clkbuf_1 _15857_ (.A(_02806_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _15858_ (.A0(net945),
    .A1(_02654_),
    .S(_02805_),
    .X(_02807_));
 sky130_fd_sc_hd__clkbuf_1 _15859_ (.A(_02807_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _15860_ (.A0(net902),
    .A1(_02656_),
    .S(_02805_),
    .X(_02808_));
 sky130_fd_sc_hd__clkbuf_1 _15861_ (.A(_02808_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _15862_ (.A0(net1325),
    .A1(_02658_),
    .S(_02805_),
    .X(_02809_));
 sky130_fd_sc_hd__clkbuf_1 _15863_ (.A(_02809_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _15864_ (.A0(net455),
    .A1(_02660_),
    .S(_02805_),
    .X(_02810_));
 sky130_fd_sc_hd__clkbuf_1 _15865_ (.A(_02810_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _15866_ (.A0(net327),
    .A1(_02662_),
    .S(_02805_),
    .X(_02811_));
 sky130_fd_sc_hd__clkbuf_1 _15867_ (.A(_02811_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _15868_ (.A0(net873),
    .A1(_02664_),
    .S(_02805_),
    .X(_02812_));
 sky130_fd_sc_hd__clkbuf_1 _15869_ (.A(_02812_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _15870_ (.A0(net892),
    .A1(_02666_),
    .S(_02805_),
    .X(_02813_));
 sky130_fd_sc_hd__clkbuf_1 _15871_ (.A(_02813_),
    .X(_00966_));
 sky130_fd_sc_hd__clkbuf_8 _15872_ (.A(_02327_),
    .X(_02814_));
 sky130_fd_sc_hd__and3_1 _15873_ (.A(_02750_),
    .B(_02297_),
    .C(_02718_),
    .X(_02815_));
 sky130_fd_sc_hd__buf_4 _15874_ (.A(_02815_),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_1 _15875_ (.A0(net513),
    .A1(_02814_),
    .S(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__clkbuf_1 _15876_ (.A(_02817_),
    .X(_00967_));
 sky130_fd_sc_hd__buf_8 _15877_ (.A(_02332_),
    .X(_02818_));
 sky130_fd_sc_hd__mux2_1 _15878_ (.A0(net1132),
    .A1(_02818_),
    .S(_02816_),
    .X(_02819_));
 sky130_fd_sc_hd__clkbuf_1 _15879_ (.A(_02819_),
    .X(_00968_));
 sky130_fd_sc_hd__buf_6 _15880_ (.A(_02335_),
    .X(_02820_));
 sky130_fd_sc_hd__mux2_1 _15881_ (.A0(net650),
    .A1(_02820_),
    .S(_02816_),
    .X(_02821_));
 sky130_fd_sc_hd__clkbuf_1 _15882_ (.A(_02821_),
    .X(_00969_));
 sky130_fd_sc_hd__clkbuf_8 _15883_ (.A(_02338_),
    .X(_02822_));
 sky130_fd_sc_hd__mux2_1 _15884_ (.A0(net486),
    .A1(_02822_),
    .S(_02816_),
    .X(_02823_));
 sky130_fd_sc_hd__clkbuf_1 _15885_ (.A(_02823_),
    .X(_00970_));
 sky130_fd_sc_hd__clkbuf_8 _15886_ (.A(_02341_),
    .X(_02824_));
 sky130_fd_sc_hd__mux2_1 _15887_ (.A0(net388),
    .A1(_02824_),
    .S(_02816_),
    .X(_02825_));
 sky130_fd_sc_hd__clkbuf_1 _15888_ (.A(_02825_),
    .X(_00971_));
 sky130_fd_sc_hd__buf_6 _15889_ (.A(_02344_),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _15890_ (.A0(net419),
    .A1(_02826_),
    .S(_02816_),
    .X(_02827_));
 sky130_fd_sc_hd__clkbuf_1 _15891_ (.A(_02827_),
    .X(_00972_));
 sky130_fd_sc_hd__buf_12 _15892_ (.A(_02347_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _15893_ (.A0(net1852),
    .A1(_02828_),
    .S(_02816_),
    .X(_02829_));
 sky130_fd_sc_hd__clkbuf_1 _15894_ (.A(_02829_),
    .X(_00973_));
 sky130_fd_sc_hd__buf_6 _15895_ (.A(_02350_),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_1 _15896_ (.A0(net697),
    .A1(_02830_),
    .S(_02816_),
    .X(_02831_));
 sky130_fd_sc_hd__clkbuf_1 _15897_ (.A(_02831_),
    .X(_00974_));
 sky130_fd_sc_hd__and3_1 _15898_ (.A(_02750_),
    .B(_08839_),
    .C(_02718_),
    .X(_02832_));
 sky130_fd_sc_hd__buf_8 _15899_ (.A(_02832_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _15900_ (.A0(net479),
    .A1(_02814_),
    .S(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__clkbuf_1 _15901_ (.A(_02834_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _15902_ (.A0(net329),
    .A1(_02818_),
    .S(_02833_),
    .X(_02835_));
 sky130_fd_sc_hd__clkbuf_1 _15903_ (.A(_02835_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _15904_ (.A0(net351),
    .A1(_02820_),
    .S(_02833_),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _15905_ (.A(_02836_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _15906_ (.A0(net854),
    .A1(_02822_),
    .S(_02833_),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_1 _15907_ (.A(_02837_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _15908_ (.A0(net993),
    .A1(_02824_),
    .S(_02833_),
    .X(_02838_));
 sky130_fd_sc_hd__clkbuf_1 _15909_ (.A(_02838_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _15910_ (.A0(net901),
    .A1(_02826_),
    .S(_02833_),
    .X(_02839_));
 sky130_fd_sc_hd__clkbuf_1 _15911_ (.A(_02839_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _15912_ (.A0(net1071),
    .A1(_02828_),
    .S(_02833_),
    .X(_02840_));
 sky130_fd_sc_hd__clkbuf_1 _15913_ (.A(_02840_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _15914_ (.A0(net963),
    .A1(_02830_),
    .S(_02833_),
    .X(_02841_));
 sky130_fd_sc_hd__clkbuf_1 _15915_ (.A(_02841_),
    .X(_00982_));
 sky130_fd_sc_hd__nand2_8 _15916_ (.A(_05985_),
    .B(_02552_),
    .Y(_02842_));
 sky130_fd_sc_hd__mux2_1 _15917_ (.A0(_02749_),
    .A1(net1950),
    .S(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__clkbuf_1 _15918_ (.A(_02843_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _15919_ (.A0(_02753_),
    .A1(\cur_mb_mem[104][1] ),
    .S(_02842_),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _15920_ (.A(_02844_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _15921_ (.A0(_02755_),
    .A1(net1944),
    .S(_02842_),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _15922_ (.A(_02845_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _15923_ (.A0(_02757_),
    .A1(\cur_mb_mem[104][3] ),
    .S(_02842_),
    .X(_02846_));
 sky130_fd_sc_hd__clkbuf_1 _15924_ (.A(_02846_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _15925_ (.A0(_02759_),
    .A1(\cur_mb_mem[104][4] ),
    .S(_02842_),
    .X(_02847_));
 sky130_fd_sc_hd__clkbuf_1 _15926_ (.A(_02847_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _15927_ (.A0(_02761_),
    .A1(\cur_mb_mem[104][5] ),
    .S(_02842_),
    .X(_02848_));
 sky130_fd_sc_hd__clkbuf_1 _15928_ (.A(_02848_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _15929_ (.A0(_02763_),
    .A1(net1742),
    .S(_02842_),
    .X(_02849_));
 sky130_fd_sc_hd__clkbuf_1 _15930_ (.A(_02849_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _15931_ (.A0(_02765_),
    .A1(\cur_mb_mem[104][7] ),
    .S(_02842_),
    .X(_02850_));
 sky130_fd_sc_hd__clkbuf_1 _15932_ (.A(_02850_),
    .X(_00990_));
 sky130_fd_sc_hd__and3_1 _15933_ (.A(_08978_),
    .B(_02750_),
    .C(_02718_),
    .X(_02851_));
 sky130_fd_sc_hd__buf_8 _15934_ (.A(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__mux2_1 _15935_ (.A0(net532),
    .A1(_02814_),
    .S(_02852_),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_1 _15936_ (.A(_02853_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _15937_ (.A0(net630),
    .A1(_02818_),
    .S(_02852_),
    .X(_02854_));
 sky130_fd_sc_hd__clkbuf_1 _15938_ (.A(_02854_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _15939_ (.A0(net1717),
    .A1(_02820_),
    .S(_02852_),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_1 _15940_ (.A(_02855_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _15941_ (.A0(net328),
    .A1(_02822_),
    .S(_02852_),
    .X(_02856_));
 sky130_fd_sc_hd__clkbuf_1 _15942_ (.A(_02856_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _15943_ (.A0(net349),
    .A1(_02824_),
    .S(_02852_),
    .X(_02857_));
 sky130_fd_sc_hd__clkbuf_1 _15944_ (.A(_02857_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _15945_ (.A0(net515),
    .A1(_02826_),
    .S(_02852_),
    .X(_02858_));
 sky130_fd_sc_hd__clkbuf_1 _15946_ (.A(_02858_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _15947_ (.A0(net1691),
    .A1(_02828_),
    .S(_02852_),
    .X(_02859_));
 sky130_fd_sc_hd__clkbuf_1 _15948_ (.A(_02859_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _15949_ (.A0(net1051),
    .A1(_02830_),
    .S(_02852_),
    .X(_02860_));
 sky130_fd_sc_hd__clkbuf_1 _15950_ (.A(_02860_),
    .X(_00998_));
 sky130_fd_sc_hd__and3_1 _15951_ (.A(_02353_),
    .B(_02750_),
    .C(_02718_),
    .X(_02861_));
 sky130_fd_sc_hd__clkbuf_8 _15952_ (.A(_02861_),
    .X(_02862_));
 sky130_fd_sc_hd__mux2_1 _15953_ (.A0(net464),
    .A1(_02814_),
    .S(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__clkbuf_1 _15954_ (.A(_02863_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _15955_ (.A0(net574),
    .A1(_02818_),
    .S(_02862_),
    .X(_02864_));
 sky130_fd_sc_hd__clkbuf_1 _15956_ (.A(_02864_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _15957_ (.A0(net482),
    .A1(_02820_),
    .S(_02862_),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_1 _15958_ (.A(_02865_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _15959_ (.A0(net499),
    .A1(_02822_),
    .S(_02862_),
    .X(_02866_));
 sky130_fd_sc_hd__clkbuf_1 _15960_ (.A(_02866_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _15961_ (.A0(net357),
    .A1(_02824_),
    .S(_02862_),
    .X(_02867_));
 sky130_fd_sc_hd__clkbuf_1 _15962_ (.A(_02867_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _15963_ (.A0(net958),
    .A1(_02826_),
    .S(_02862_),
    .X(_02868_));
 sky130_fd_sc_hd__clkbuf_1 _15964_ (.A(_02868_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _15965_ (.A0(net1437),
    .A1(_02828_),
    .S(_02862_),
    .X(_02869_));
 sky130_fd_sc_hd__clkbuf_1 _15966_ (.A(_02869_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _15967_ (.A0(net789),
    .A1(_02830_),
    .S(_02862_),
    .X(_02870_));
 sky130_fd_sc_hd__clkbuf_1 _15968_ (.A(_02870_),
    .X(_01006_));
 sky130_fd_sc_hd__and3_1 _15969_ (.A(_02526_),
    .B(_02750_),
    .C(_02718_),
    .X(_02871_));
 sky130_fd_sc_hd__clkbuf_8 _15970_ (.A(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_1 _15971_ (.A0(net1049),
    .A1(_02814_),
    .S(_02872_),
    .X(_02873_));
 sky130_fd_sc_hd__clkbuf_1 _15972_ (.A(_02873_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _15973_ (.A0(net462),
    .A1(_02818_),
    .S(_02872_),
    .X(_02874_));
 sky130_fd_sc_hd__clkbuf_1 _15974_ (.A(_02874_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _15975_ (.A0(net439),
    .A1(_02820_),
    .S(_02872_),
    .X(_02875_));
 sky130_fd_sc_hd__clkbuf_1 _15976_ (.A(_02875_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _15977_ (.A0(net548),
    .A1(_02822_),
    .S(_02872_),
    .X(_02876_));
 sky130_fd_sc_hd__clkbuf_1 _15978_ (.A(_02876_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _15979_ (.A0(net580),
    .A1(_02824_),
    .S(_02872_),
    .X(_02877_));
 sky130_fd_sc_hd__clkbuf_1 _15980_ (.A(_02877_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _15981_ (.A0(net644),
    .A1(_02826_),
    .S(_02872_),
    .X(_02878_));
 sky130_fd_sc_hd__clkbuf_1 _15982_ (.A(_02878_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _15983_ (.A0(net918),
    .A1(_02828_),
    .S(_02872_),
    .X(_02879_));
 sky130_fd_sc_hd__clkbuf_1 _15984_ (.A(_02879_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _15985_ (.A0(net1904),
    .A1(_02830_),
    .S(_02872_),
    .X(_02880_));
 sky130_fd_sc_hd__clkbuf_1 _15986_ (.A(_02880_),
    .X(_01014_));
 sky130_fd_sc_hd__clkbuf_4 _15987_ (.A(_08900_),
    .X(_02881_));
 sky130_fd_sc_hd__and3_1 _15988_ (.A(_02374_),
    .B(_06299_),
    .C(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__buf_12 _15989_ (.A(_02882_),
    .X(_02883_));
 sky130_fd_sc_hd__mux2_1 _15990_ (.A0(net1835),
    .A1(_02814_),
    .S(_02883_),
    .X(_02884_));
 sky130_fd_sc_hd__clkbuf_1 _15991_ (.A(_02884_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _15992_ (.A0(net316),
    .A1(_02818_),
    .S(_02883_),
    .X(_02885_));
 sky130_fd_sc_hd__clkbuf_1 _15993_ (.A(_02885_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _15994_ (.A0(net1863),
    .A1(_02820_),
    .S(_02883_),
    .X(_02886_));
 sky130_fd_sc_hd__clkbuf_1 _15995_ (.A(_02886_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _15996_ (.A0(net1849),
    .A1(_02822_),
    .S(_02883_),
    .X(_02887_));
 sky130_fd_sc_hd__clkbuf_1 _15997_ (.A(_02887_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _15998_ (.A0(net837),
    .A1(_02824_),
    .S(_02883_),
    .X(_02888_));
 sky130_fd_sc_hd__clkbuf_1 _15999_ (.A(_02888_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _16000_ (.A0(net1207),
    .A1(_02826_),
    .S(_02883_),
    .X(_02889_));
 sky130_fd_sc_hd__clkbuf_1 _16001_ (.A(_02889_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _16002_ (.A0(net1550),
    .A1(_02828_),
    .S(_02883_),
    .X(_02890_));
 sky130_fd_sc_hd__clkbuf_1 _16003_ (.A(_02890_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _16004_ (.A0(net1387),
    .A1(_02830_),
    .S(_02883_),
    .X(_02891_));
 sky130_fd_sc_hd__clkbuf_1 _16005_ (.A(_02891_),
    .X(_01022_));
 sky130_fd_sc_hd__and3_1 _16006_ (.A(_02750_),
    .B(_05961_),
    .C(_02881_),
    .X(_02892_));
 sky130_fd_sc_hd__buf_4 _16007_ (.A(_02892_),
    .X(_02893_));
 sky130_fd_sc_hd__mux2_1 _16008_ (.A0(net638),
    .A1(_02814_),
    .S(_02893_),
    .X(_02894_));
 sky130_fd_sc_hd__clkbuf_1 _16009_ (.A(_02894_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _16010_ (.A0(net456),
    .A1(_02818_),
    .S(_02893_),
    .X(_02895_));
 sky130_fd_sc_hd__clkbuf_1 _16011_ (.A(_02895_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _16012_ (.A0(net344),
    .A1(_02820_),
    .S(_02893_),
    .X(_02896_));
 sky130_fd_sc_hd__clkbuf_1 _16013_ (.A(_02896_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _16014_ (.A0(net402),
    .A1(_02822_),
    .S(_02893_),
    .X(_02897_));
 sky130_fd_sc_hd__clkbuf_1 _16015_ (.A(_02897_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _16016_ (.A0(net330),
    .A1(_02824_),
    .S(_02893_),
    .X(_02898_));
 sky130_fd_sc_hd__clkbuf_1 _16017_ (.A(_02898_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _16018_ (.A0(net672),
    .A1(_02826_),
    .S(_02893_),
    .X(_02899_));
 sky130_fd_sc_hd__clkbuf_1 _16019_ (.A(_02899_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _16020_ (.A0(net1082),
    .A1(_02828_),
    .S(_02893_),
    .X(_02900_));
 sky130_fd_sc_hd__clkbuf_1 _16021_ (.A(_02900_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _16022_ (.A0(net859),
    .A1(_02830_),
    .S(_02893_),
    .X(_02901_));
 sky130_fd_sc_hd__clkbuf_1 _16023_ (.A(_02901_),
    .X(_01030_));
 sky130_fd_sc_hd__and3_1 _16024_ (.A(_02750_),
    .B(_09036_),
    .C(_02881_),
    .X(_02902_));
 sky130_fd_sc_hd__clkbuf_8 _16025_ (.A(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__mux2_1 _16026_ (.A0(net1519),
    .A1(_02814_),
    .S(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__clkbuf_1 _16027_ (.A(_02904_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _16028_ (.A0(net824),
    .A1(_02818_),
    .S(_02903_),
    .X(_02905_));
 sky130_fd_sc_hd__clkbuf_1 _16029_ (.A(_02905_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _16030_ (.A0(net1084),
    .A1(_02820_),
    .S(_02903_),
    .X(_02906_));
 sky130_fd_sc_hd__clkbuf_1 _16031_ (.A(_02906_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _16032_ (.A0(net785),
    .A1(_02822_),
    .S(_02903_),
    .X(_02907_));
 sky130_fd_sc_hd__clkbuf_1 _16033_ (.A(_02907_),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_1 _16034_ (.A0(net885),
    .A1(_02824_),
    .S(_02903_),
    .X(_02908_));
 sky130_fd_sc_hd__clkbuf_1 _16035_ (.A(_02908_),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _16036_ (.A0(net1440),
    .A1(_02826_),
    .S(_02903_),
    .X(_02909_));
 sky130_fd_sc_hd__clkbuf_1 _16037_ (.A(_02909_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _16038_ (.A0(net1345),
    .A1(_02828_),
    .S(_02903_),
    .X(_02910_));
 sky130_fd_sc_hd__clkbuf_1 _16039_ (.A(_02910_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _16040_ (.A0(net813),
    .A1(_02830_),
    .S(_02903_),
    .X(_02911_));
 sky130_fd_sc_hd__clkbuf_1 _16041_ (.A(_02911_),
    .X(_01038_));
 sky130_fd_sc_hd__and3_1 _16042_ (.A(_02406_),
    .B(_06299_),
    .C(_02881_),
    .X(_02912_));
 sky130_fd_sc_hd__clkbuf_16 _16043_ (.A(_02912_),
    .X(_02913_));
 sky130_fd_sc_hd__mux2_1 _16044_ (.A0(net379),
    .A1(_02814_),
    .S(_02913_),
    .X(_02914_));
 sky130_fd_sc_hd__clkbuf_1 _16045_ (.A(_02914_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _16046_ (.A0(net1680),
    .A1(_02818_),
    .S(_02913_),
    .X(_02915_));
 sky130_fd_sc_hd__clkbuf_1 _16047_ (.A(_02915_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _16048_ (.A0(net318),
    .A1(_02820_),
    .S(_02913_),
    .X(_02916_));
 sky130_fd_sc_hd__clkbuf_1 _16049_ (.A(_02916_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _16050_ (.A0(net334),
    .A1(_02822_),
    .S(_02913_),
    .X(_02917_));
 sky130_fd_sc_hd__clkbuf_1 _16051_ (.A(_02917_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _16052_ (.A0(net786),
    .A1(_02824_),
    .S(_02913_),
    .X(_02918_));
 sky130_fd_sc_hd__clkbuf_1 _16053_ (.A(_02918_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _16054_ (.A0(net920),
    .A1(_02826_),
    .S(_02913_),
    .X(_02919_));
 sky130_fd_sc_hd__clkbuf_1 _16055_ (.A(_02919_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _16056_ (.A0(net818),
    .A1(_02828_),
    .S(_02913_),
    .X(_02920_));
 sky130_fd_sc_hd__clkbuf_1 _16057_ (.A(_02920_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _16058_ (.A0(net1128),
    .A1(_02830_),
    .S(_02913_),
    .X(_02921_));
 sky130_fd_sc_hd__clkbuf_1 _16059_ (.A(_02921_),
    .X(_01046_));
 sky130_fd_sc_hd__clkbuf_4 _16060_ (.A(_06119_),
    .X(_02922_));
 sky130_fd_sc_hd__nand2_4 _16061_ (.A(_02922_),
    .B(_08883_),
    .Y(_02923_));
 sky130_fd_sc_hd__mux2_1 _16062_ (.A0(_02749_),
    .A1(net1747),
    .S(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__clkbuf_1 _16063_ (.A(_02924_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _16064_ (.A0(_02753_),
    .A1(\cur_mb_mem[112][1] ),
    .S(_02923_),
    .X(_02925_));
 sky130_fd_sc_hd__clkbuf_1 _16065_ (.A(_02925_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _16066_ (.A0(_02755_),
    .A1(net1801),
    .S(_02923_),
    .X(_02926_));
 sky130_fd_sc_hd__clkbuf_1 _16067_ (.A(_02926_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _16068_ (.A0(_02757_),
    .A1(\cur_mb_mem[112][3] ),
    .S(_02923_),
    .X(_02927_));
 sky130_fd_sc_hd__clkbuf_1 _16069_ (.A(_02927_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _16070_ (.A0(_02759_),
    .A1(net1477),
    .S(_02923_),
    .X(_02928_));
 sky130_fd_sc_hd__clkbuf_1 _16071_ (.A(_02928_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _16072_ (.A0(_02761_),
    .A1(net1667),
    .S(_02923_),
    .X(_02929_));
 sky130_fd_sc_hd__clkbuf_1 _16073_ (.A(_02929_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _16074_ (.A0(_02763_),
    .A1(\cur_mb_mem[112][6] ),
    .S(_02923_),
    .X(_02930_));
 sky130_fd_sc_hd__clkbuf_1 _16075_ (.A(_02930_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _16076_ (.A0(_02765_),
    .A1(\cur_mb_mem[112][7] ),
    .S(_02923_),
    .X(_02931_));
 sky130_fd_sc_hd__clkbuf_1 _16077_ (.A(_02931_),
    .X(_01054_));
 sky130_fd_sc_hd__nand3_4 _16078_ (.A(_02922_),
    .B(_05994_),
    .C(_08901_),
    .Y(_02932_));
 sky130_fd_sc_hd__mux2_1 _16079_ (.A0(_02749_),
    .A1(\cur_mb_mem[113][0] ),
    .S(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__clkbuf_1 _16080_ (.A(_02933_),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _16081_ (.A0(_02753_),
    .A1(\cur_mb_mem[113][1] ),
    .S(_02932_),
    .X(_02934_));
 sky130_fd_sc_hd__clkbuf_1 _16082_ (.A(_02934_),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _16083_ (.A0(_02755_),
    .A1(net1564),
    .S(_02932_),
    .X(_02935_));
 sky130_fd_sc_hd__clkbuf_1 _16084_ (.A(_02935_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _16085_ (.A0(_02757_),
    .A1(\cur_mb_mem[113][3] ),
    .S(_02932_),
    .X(_02936_));
 sky130_fd_sc_hd__clkbuf_1 _16086_ (.A(_02936_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _16087_ (.A0(_02759_),
    .A1(net1590),
    .S(_02932_),
    .X(_02937_));
 sky130_fd_sc_hd__clkbuf_1 _16088_ (.A(_02937_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _16089_ (.A0(_02761_),
    .A1(net1496),
    .S(_02932_),
    .X(_02938_));
 sky130_fd_sc_hd__clkbuf_1 _16090_ (.A(_02938_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _16091_ (.A0(_02763_),
    .A1(\cur_mb_mem[113][6] ),
    .S(_02932_),
    .X(_02939_));
 sky130_fd_sc_hd__clkbuf_1 _16092_ (.A(_02939_),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _16093_ (.A0(_02765_),
    .A1(\cur_mb_mem[113][7] ),
    .S(_02932_),
    .X(_02940_));
 sky130_fd_sc_hd__clkbuf_1 _16094_ (.A(_02940_),
    .X(_01062_));
 sky130_fd_sc_hd__nand2_8 _16095_ (.A(_06280_),
    .B(_02552_),
    .Y(_02941_));
 sky130_fd_sc_hd__mux2_1 _16096_ (.A0(_02749_),
    .A1(\cur_mb_mem[114][0] ),
    .S(_02941_),
    .X(_02942_));
 sky130_fd_sc_hd__clkbuf_1 _16097_ (.A(_02942_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _16098_ (.A0(_02753_),
    .A1(\cur_mb_mem[114][1] ),
    .S(_02941_),
    .X(_02943_));
 sky130_fd_sc_hd__clkbuf_1 _16099_ (.A(_02943_),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _16100_ (.A0(_02755_),
    .A1(net1773),
    .S(_02941_),
    .X(_02944_));
 sky130_fd_sc_hd__clkbuf_1 _16101_ (.A(_02944_),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _16102_ (.A0(_02757_),
    .A1(\cur_mb_mem[114][3] ),
    .S(_02941_),
    .X(_02945_));
 sky130_fd_sc_hd__clkbuf_1 _16103_ (.A(_02945_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _16104_ (.A0(_02759_),
    .A1(net1731),
    .S(_02941_),
    .X(_02946_));
 sky130_fd_sc_hd__clkbuf_1 _16105_ (.A(_02946_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _16106_ (.A0(_02761_),
    .A1(net1724),
    .S(_02941_),
    .X(_02947_));
 sky130_fd_sc_hd__clkbuf_1 _16107_ (.A(_02947_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _16108_ (.A0(_02763_),
    .A1(\cur_mb_mem[114][6] ),
    .S(_02941_),
    .X(_02948_));
 sky130_fd_sc_hd__clkbuf_1 _16109_ (.A(_02948_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _16110_ (.A0(_02765_),
    .A1(\cur_mb_mem[114][7] ),
    .S(_02941_),
    .X(_02949_));
 sky130_fd_sc_hd__clkbuf_1 _16111_ (.A(_02949_),
    .X(_01070_));
 sky130_fd_sc_hd__and3_1 _16112_ (.A(_02266_),
    .B(_02922_),
    .C(_02881_),
    .X(_02950_));
 sky130_fd_sc_hd__buf_8 _16113_ (.A(_02950_),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_1 _16114_ (.A0(net1726),
    .A1(_02814_),
    .S(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__clkbuf_1 _16115_ (.A(_02952_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _16116_ (.A0(net473),
    .A1(_02818_),
    .S(_02951_),
    .X(_02953_));
 sky130_fd_sc_hd__clkbuf_1 _16117_ (.A(_02953_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _16118_ (.A0(net1675),
    .A1(_02820_),
    .S(_02951_),
    .X(_02954_));
 sky130_fd_sc_hd__clkbuf_1 _16119_ (.A(_02954_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _16120_ (.A0(net480),
    .A1(_02822_),
    .S(_02951_),
    .X(_02955_));
 sky130_fd_sc_hd__clkbuf_1 _16121_ (.A(_02955_),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _16122_ (.A0(net414),
    .A1(_02824_),
    .S(_02951_),
    .X(_02956_));
 sky130_fd_sc_hd__clkbuf_1 _16123_ (.A(_02956_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _16124_ (.A0(net366),
    .A1(_02826_),
    .S(_02951_),
    .X(_02957_));
 sky130_fd_sc_hd__clkbuf_1 _16125_ (.A(_02957_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _16126_ (.A0(net1596),
    .A1(_02828_),
    .S(_02951_),
    .X(_02958_));
 sky130_fd_sc_hd__clkbuf_1 _16127_ (.A(_02958_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _16128_ (.A0(net444),
    .A1(_02830_),
    .S(_02951_),
    .X(_02959_));
 sky130_fd_sc_hd__clkbuf_1 _16129_ (.A(_02959_),
    .X(_01078_));
 sky130_fd_sc_hd__nand2_4 _16130_ (.A(_06239_),
    .B(_02552_),
    .Y(_02960_));
 sky130_fd_sc_hd__mux2_1 _16131_ (.A0(_02749_),
    .A1(\cur_mb_mem[116][0] ),
    .S(_02960_),
    .X(_02961_));
 sky130_fd_sc_hd__clkbuf_1 _16132_ (.A(_02961_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _16133_ (.A0(_02753_),
    .A1(\cur_mb_mem[116][1] ),
    .S(_02960_),
    .X(_02962_));
 sky130_fd_sc_hd__clkbuf_1 _16134_ (.A(_02962_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _16135_ (.A0(_02755_),
    .A1(net1983),
    .S(_02960_),
    .X(_02963_));
 sky130_fd_sc_hd__clkbuf_1 _16136_ (.A(_02963_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _16137_ (.A0(_02757_),
    .A1(\cur_mb_mem[116][3] ),
    .S(_02960_),
    .X(_02964_));
 sky130_fd_sc_hd__clkbuf_1 _16138_ (.A(_02964_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _16139_ (.A0(_02759_),
    .A1(net1453),
    .S(_02960_),
    .X(_02965_));
 sky130_fd_sc_hd__clkbuf_1 _16140_ (.A(_02965_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _16141_ (.A0(_02761_),
    .A1(net1421),
    .S(_02960_),
    .X(_02966_));
 sky130_fd_sc_hd__clkbuf_1 _16142_ (.A(_02966_),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _16143_ (.A0(_02763_),
    .A1(\cur_mb_mem[116][6] ),
    .S(_02960_),
    .X(_02967_));
 sky130_fd_sc_hd__clkbuf_1 _16144_ (.A(_02967_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _16145_ (.A0(_02765_),
    .A1(\cur_mb_mem[116][7] ),
    .S(_02960_),
    .X(_02968_));
 sky130_fd_sc_hd__clkbuf_1 _16146_ (.A(_02968_),
    .X(_01086_));
 sky130_fd_sc_hd__buf_8 _16147_ (.A(_02327_),
    .X(_02969_));
 sky130_fd_sc_hd__and3_1 _16148_ (.A(_02922_),
    .B(_02286_),
    .C(_02881_),
    .X(_02970_));
 sky130_fd_sc_hd__buf_4 _16149_ (.A(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__mux2_1 _16150_ (.A0(net386),
    .A1(_02969_),
    .S(_02971_),
    .X(_02972_));
 sky130_fd_sc_hd__clkbuf_1 _16151_ (.A(_02972_),
    .X(_01087_));
 sky130_fd_sc_hd__buf_8 _16152_ (.A(_02332_),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_1 _16153_ (.A0(\cur_mb_mem[117][1] ),
    .A1(_02973_),
    .S(_02971_),
    .X(_02974_));
 sky130_fd_sc_hd__clkbuf_1 _16154_ (.A(_02974_),
    .X(_01088_));
 sky130_fd_sc_hd__buf_8 _16155_ (.A(_02335_),
    .X(_02975_));
 sky130_fd_sc_hd__mux2_1 _16156_ (.A0(net688),
    .A1(_02975_),
    .S(_02971_),
    .X(_02976_));
 sky130_fd_sc_hd__clkbuf_1 _16157_ (.A(_02976_),
    .X(_01089_));
 sky130_fd_sc_hd__buf_8 _16158_ (.A(_02338_),
    .X(_02977_));
 sky130_fd_sc_hd__mux2_1 _16159_ (.A0(net341),
    .A1(_02977_),
    .S(_02971_),
    .X(_02978_));
 sky130_fd_sc_hd__clkbuf_1 _16160_ (.A(_02978_),
    .X(_01090_));
 sky130_fd_sc_hd__buf_6 _16161_ (.A(_02341_),
    .X(_02979_));
 sky130_fd_sc_hd__mux2_1 _16162_ (.A0(net1621),
    .A1(_02979_),
    .S(_02971_),
    .X(_02980_));
 sky130_fd_sc_hd__clkbuf_1 _16163_ (.A(_02980_),
    .X(_01091_));
 sky130_fd_sc_hd__buf_6 _16164_ (.A(_02344_),
    .X(_02981_));
 sky130_fd_sc_hd__mux2_1 _16165_ (.A0(net1572),
    .A1(_02981_),
    .S(_02971_),
    .X(_02982_));
 sky130_fd_sc_hd__clkbuf_1 _16166_ (.A(_02982_),
    .X(_01092_));
 sky130_fd_sc_hd__buf_6 _16167_ (.A(_02347_),
    .X(_02983_));
 sky130_fd_sc_hd__mux2_1 _16168_ (.A0(\cur_mb_mem[117][6] ),
    .A1(_02983_),
    .S(_02971_),
    .X(_02984_));
 sky130_fd_sc_hd__clkbuf_1 _16169_ (.A(_02984_),
    .X(_01093_));
 sky130_fd_sc_hd__buf_8 _16170_ (.A(_02350_),
    .X(_02985_));
 sky130_fd_sc_hd__mux2_1 _16171_ (.A0(\cur_mb_mem[117][7] ),
    .A1(_02985_),
    .S(_02971_),
    .X(_02986_));
 sky130_fd_sc_hd__clkbuf_1 _16172_ (.A(_02986_),
    .X(_01094_));
 sky130_fd_sc_hd__and3_1 _16173_ (.A(_02922_),
    .B(_02297_),
    .C(_02881_),
    .X(_02987_));
 sky130_fd_sc_hd__buf_6 _16174_ (.A(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _16175_ (.A0(net1399),
    .A1(_02969_),
    .S(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__clkbuf_1 _16176_ (.A(_02989_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _16177_ (.A0(net1154),
    .A1(_02973_),
    .S(_02988_),
    .X(_02990_));
 sky130_fd_sc_hd__clkbuf_1 _16178_ (.A(_02990_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _16179_ (.A0(net1673),
    .A1(_02975_),
    .S(_02988_),
    .X(_02991_));
 sky130_fd_sc_hd__clkbuf_1 _16180_ (.A(_02991_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _16181_ (.A0(net988),
    .A1(_02977_),
    .S(_02988_),
    .X(_02992_));
 sky130_fd_sc_hd__clkbuf_1 _16182_ (.A(_02992_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _16183_ (.A0(net1034),
    .A1(_02979_),
    .S(_02988_),
    .X(_02993_));
 sky130_fd_sc_hd__clkbuf_1 _16184_ (.A(_02993_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _16185_ (.A0(net1095),
    .A1(_02981_),
    .S(_02988_),
    .X(_02994_));
 sky130_fd_sc_hd__clkbuf_1 _16186_ (.A(_02994_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _16187_ (.A0(net1011),
    .A1(_02983_),
    .S(_02988_),
    .X(_02995_));
 sky130_fd_sc_hd__clkbuf_1 _16188_ (.A(_02995_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _16189_ (.A0(net1293),
    .A1(_02985_),
    .S(_02988_),
    .X(_02996_));
 sky130_fd_sc_hd__clkbuf_1 _16190_ (.A(_02996_),
    .X(_01102_));
 sky130_fd_sc_hd__and3_1 _16191_ (.A(_02922_),
    .B(_08839_),
    .C(_02881_),
    .X(_02997_));
 sky130_fd_sc_hd__buf_6 _16192_ (.A(_02997_),
    .X(_02998_));
 sky130_fd_sc_hd__mux2_1 _16193_ (.A0(net422),
    .A1(_02969_),
    .S(_02998_),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_1 _16194_ (.A(_02999_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _16195_ (.A0(net543),
    .A1(_02973_),
    .S(_02998_),
    .X(_03000_));
 sky130_fd_sc_hd__clkbuf_1 _16196_ (.A(_03000_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _16197_ (.A0(net435),
    .A1(_02975_),
    .S(_02998_),
    .X(_03001_));
 sky130_fd_sc_hd__clkbuf_1 _16198_ (.A(_03001_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _16199_ (.A0(net1000),
    .A1(_02977_),
    .S(_02998_),
    .X(_03002_));
 sky130_fd_sc_hd__clkbuf_1 _16200_ (.A(_03002_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _16201_ (.A0(net1687),
    .A1(_02979_),
    .S(_02998_),
    .X(_03003_));
 sky130_fd_sc_hd__clkbuf_1 _16202_ (.A(_03003_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _16203_ (.A0(net1779),
    .A1(_02981_),
    .S(_02998_),
    .X(_03004_));
 sky130_fd_sc_hd__clkbuf_1 _16204_ (.A(_03004_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _16205_ (.A0(net1197),
    .A1(_02983_),
    .S(_02998_),
    .X(_03005_));
 sky130_fd_sc_hd__clkbuf_1 _16206_ (.A(_03005_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _16207_ (.A0(net742),
    .A1(_02985_),
    .S(_02998_),
    .X(_03006_));
 sky130_fd_sc_hd__clkbuf_1 _16208_ (.A(_03006_),
    .X(_01110_));
 sky130_fd_sc_hd__nand2_8 _16209_ (.A(_06432_),
    .B(_02552_),
    .Y(_03007_));
 sky130_fd_sc_hd__mux2_1 _16210_ (.A0(_02749_),
    .A1(net1671),
    .S(_03007_),
    .X(_03008_));
 sky130_fd_sc_hd__clkbuf_1 _16211_ (.A(_03008_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _16212_ (.A0(_02753_),
    .A1(net1793),
    .S(_03007_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_1 _16213_ (.A(_03009_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _16214_ (.A0(_02755_),
    .A1(net1825),
    .S(_03007_),
    .X(_03010_));
 sky130_fd_sc_hd__clkbuf_1 _16215_ (.A(_03010_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _16216_ (.A0(_02757_),
    .A1(net1847),
    .S(_03007_),
    .X(_03011_));
 sky130_fd_sc_hd__clkbuf_1 _16217_ (.A(_03011_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _16218_ (.A0(_02759_),
    .A1(net1897),
    .S(_03007_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_1 _16219_ (.A(_03012_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _16220_ (.A0(_02761_),
    .A1(net1853),
    .S(_03007_),
    .X(_03013_));
 sky130_fd_sc_hd__clkbuf_1 _16221_ (.A(_03013_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _16222_ (.A0(_02763_),
    .A1(\cur_mb_mem[120][6] ),
    .S(_03007_),
    .X(_03014_));
 sky130_fd_sc_hd__clkbuf_1 _16223_ (.A(_03014_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _16224_ (.A0(_02765_),
    .A1(\cur_mb_mem[120][7] ),
    .S(_03007_),
    .X(_03015_));
 sky130_fd_sc_hd__clkbuf_1 _16225_ (.A(_03015_),
    .X(_01118_));
 sky130_fd_sc_hd__and3_1 _16226_ (.A(_08978_),
    .B(_02922_),
    .C(_02881_),
    .X(_03016_));
 sky130_fd_sc_hd__buf_4 _16227_ (.A(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__mux2_1 _16228_ (.A0(net590),
    .A1(_02969_),
    .S(_03017_),
    .X(_03018_));
 sky130_fd_sc_hd__clkbuf_1 _16229_ (.A(_03018_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _16230_ (.A0(net1058),
    .A1(_02973_),
    .S(_03017_),
    .X(_03019_));
 sky130_fd_sc_hd__clkbuf_1 _16231_ (.A(_03019_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _16232_ (.A0(net440),
    .A1(_02975_),
    .S(_03017_),
    .X(_03020_));
 sky130_fd_sc_hd__clkbuf_1 _16233_ (.A(_03020_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _16234_ (.A0(net647),
    .A1(_02977_),
    .S(_03017_),
    .X(_03021_));
 sky130_fd_sc_hd__clkbuf_1 _16235_ (.A(_03021_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _16236_ (.A0(net1118),
    .A1(_02979_),
    .S(_03017_),
    .X(_03022_));
 sky130_fd_sc_hd__clkbuf_1 _16237_ (.A(_03022_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _16238_ (.A0(net968),
    .A1(_02981_),
    .S(_03017_),
    .X(_03023_));
 sky130_fd_sc_hd__clkbuf_1 _16239_ (.A(_03023_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _16240_ (.A0(\cur_mb_mem[121][6] ),
    .A1(_02983_),
    .S(_03017_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_1 _16241_ (.A(_03024_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _16242_ (.A0(\cur_mb_mem[121][7] ),
    .A1(_02985_),
    .S(_03017_),
    .X(_03025_));
 sky130_fd_sc_hd__clkbuf_1 _16243_ (.A(_03025_),
    .X(_01126_));
 sky130_fd_sc_hd__and3_1 _16244_ (.A(_02353_),
    .B(_02922_),
    .C(_02881_),
    .X(_03026_));
 sky130_fd_sc_hd__buf_4 _16245_ (.A(_03026_),
    .X(_03027_));
 sky130_fd_sc_hd__mux2_1 _16246_ (.A0(net1261),
    .A1(_02969_),
    .S(_03027_),
    .X(_03028_));
 sky130_fd_sc_hd__clkbuf_1 _16247_ (.A(_03028_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _16248_ (.A0(\cur_mb_mem[122][1] ),
    .A1(_02973_),
    .S(_03027_),
    .X(_03029_));
 sky130_fd_sc_hd__clkbuf_1 _16249_ (.A(_03029_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _16250_ (.A0(net990),
    .A1(_02975_),
    .S(_03027_),
    .X(_03030_));
 sky130_fd_sc_hd__clkbuf_1 _16251_ (.A(_03030_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _16252_ (.A0(net658),
    .A1(_02977_),
    .S(_03027_),
    .X(_03031_));
 sky130_fd_sc_hd__clkbuf_1 _16253_ (.A(_03031_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _16254_ (.A0(net1702),
    .A1(_02979_),
    .S(_03027_),
    .X(_03032_));
 sky130_fd_sc_hd__clkbuf_1 _16255_ (.A(_03032_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _16256_ (.A0(net1712),
    .A1(_02981_),
    .S(_03027_),
    .X(_03033_));
 sky130_fd_sc_hd__clkbuf_1 _16257_ (.A(_03033_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _16258_ (.A0(\cur_mb_mem[122][6] ),
    .A1(_02983_),
    .S(_03027_),
    .X(_03034_));
 sky130_fd_sc_hd__clkbuf_1 _16259_ (.A(_03034_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _16260_ (.A0(net689),
    .A1(_02985_),
    .S(_03027_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_1 _16261_ (.A(_03035_),
    .X(_01134_));
 sky130_fd_sc_hd__buf_4 _16262_ (.A(_08900_),
    .X(_03036_));
 sky130_fd_sc_hd__and3_1 _16263_ (.A(_02526_),
    .B(_02922_),
    .C(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__buf_4 _16264_ (.A(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__mux2_1 _16265_ (.A0(net566),
    .A1(_02969_),
    .S(_03038_),
    .X(_03039_));
 sky130_fd_sc_hd__clkbuf_1 _16266_ (.A(_03039_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _16267_ (.A0(net426),
    .A1(_02973_),
    .S(_03038_),
    .X(_03040_));
 sky130_fd_sc_hd__clkbuf_1 _16268_ (.A(_03040_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _16269_ (.A0(net545),
    .A1(_02975_),
    .S(_03038_),
    .X(_03041_));
 sky130_fd_sc_hd__clkbuf_1 _16270_ (.A(_03041_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _16271_ (.A0(net605),
    .A1(_02977_),
    .S(_03038_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_1 _16272_ (.A(_03042_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _16273_ (.A0(net1975),
    .A1(_02979_),
    .S(_03038_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_1 _16274_ (.A(_03043_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _16275_ (.A0(\cur_mb_mem[123][5] ),
    .A1(_02981_),
    .S(_03038_),
    .X(_03044_));
 sky130_fd_sc_hd__clkbuf_1 _16276_ (.A(_03044_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _16277_ (.A0(net1648),
    .A1(_02983_),
    .S(_03038_),
    .X(_03045_));
 sky130_fd_sc_hd__clkbuf_1 _16278_ (.A(_03045_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _16279_ (.A0(net1218),
    .A1(_02985_),
    .S(_03038_),
    .X(_03046_));
 sky130_fd_sc_hd__clkbuf_1 _16280_ (.A(_03046_),
    .X(_01142_));
 sky130_fd_sc_hd__and3_1 _16281_ (.A(_02374_),
    .B(_06119_),
    .C(_03036_),
    .X(_03047_));
 sky130_fd_sc_hd__buf_4 _16282_ (.A(_03047_),
    .X(_03048_));
 sky130_fd_sc_hd__mux2_1 _16283_ (.A0(net1269),
    .A1(_02969_),
    .S(_03048_),
    .X(_03049_));
 sky130_fd_sc_hd__clkbuf_1 _16284_ (.A(_03049_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _16285_ (.A0(\cur_mb_mem[124][1] ),
    .A1(_02973_),
    .S(_03048_),
    .X(_03050_));
 sky130_fd_sc_hd__clkbuf_1 _16286_ (.A(_03050_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _16287_ (.A0(net1192),
    .A1(_02975_),
    .S(_03048_),
    .X(_03051_));
 sky130_fd_sc_hd__clkbuf_1 _16288_ (.A(_03051_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _16289_ (.A0(net1843),
    .A1(_02977_),
    .S(_03048_),
    .X(_03052_));
 sky130_fd_sc_hd__clkbuf_1 _16290_ (.A(_03052_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _16291_ (.A0(net1259),
    .A1(_02979_),
    .S(_03048_),
    .X(_03053_));
 sky130_fd_sc_hd__clkbuf_1 _16292_ (.A(_03053_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _16293_ (.A0(net827),
    .A1(_02981_),
    .S(_03048_),
    .X(_03054_));
 sky130_fd_sc_hd__clkbuf_1 _16294_ (.A(_03054_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _16295_ (.A0(net659),
    .A1(_02983_),
    .S(_03048_),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_1 _16296_ (.A(_03055_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _16297_ (.A0(\cur_mb_mem[124][7] ),
    .A1(_02985_),
    .S(_03048_),
    .X(_03056_));
 sky130_fd_sc_hd__clkbuf_1 _16298_ (.A(_03056_),
    .X(_01150_));
 sky130_fd_sc_hd__and3_1 _16299_ (.A(_09025_),
    .B(_06119_),
    .C(_03036_),
    .X(_03057_));
 sky130_fd_sc_hd__buf_4 _16300_ (.A(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__mux2_1 _16301_ (.A0(net1468),
    .A1(_02969_),
    .S(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__clkbuf_1 _16302_ (.A(_03059_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _16303_ (.A0(\cur_mb_mem[125][1] ),
    .A1(_02973_),
    .S(_03058_),
    .X(_03060_));
 sky130_fd_sc_hd__clkbuf_1 _16304_ (.A(_03060_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _16305_ (.A0(net549),
    .A1(_02975_),
    .S(_03058_),
    .X(_03061_));
 sky130_fd_sc_hd__clkbuf_1 _16306_ (.A(_03061_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _16307_ (.A0(net748),
    .A1(_02977_),
    .S(_03058_),
    .X(_03062_));
 sky130_fd_sc_hd__clkbuf_1 _16308_ (.A(_03062_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _16309_ (.A0(net387),
    .A1(_02979_),
    .S(_03058_),
    .X(_03063_));
 sky130_fd_sc_hd__clkbuf_1 _16310_ (.A(_03063_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _16311_ (.A0(net895),
    .A1(_02981_),
    .S(_03058_),
    .X(_03064_));
 sky130_fd_sc_hd__clkbuf_1 _16312_ (.A(_03064_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _16313_ (.A0(net849),
    .A1(_02983_),
    .S(_03058_),
    .X(_03065_));
 sky130_fd_sc_hd__clkbuf_1 _16314_ (.A(_03065_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _16315_ (.A0(\cur_mb_mem[125][7] ),
    .A1(_02985_),
    .S(_03058_),
    .X(_03066_));
 sky130_fd_sc_hd__clkbuf_1 _16316_ (.A(_03066_),
    .X(_01158_));
 sky130_fd_sc_hd__and3_1 _16317_ (.A(_02922_),
    .B(_09036_),
    .C(_03036_),
    .X(_03067_));
 sky130_fd_sc_hd__buf_6 _16318_ (.A(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__mux2_1 _16319_ (.A0(net732),
    .A1(_02969_),
    .S(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_1 _16320_ (.A(_03069_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _16321_ (.A0(net359),
    .A1(_02973_),
    .S(_03068_),
    .X(_03070_));
 sky130_fd_sc_hd__clkbuf_1 _16322_ (.A(_03070_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _16323_ (.A0(net746),
    .A1(_02975_),
    .S(_03068_),
    .X(_03071_));
 sky130_fd_sc_hd__clkbuf_1 _16324_ (.A(_03071_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _16325_ (.A0(net692),
    .A1(_02977_),
    .S(_03068_),
    .X(_03072_));
 sky130_fd_sc_hd__clkbuf_1 _16326_ (.A(_03072_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _16327_ (.A0(net1693),
    .A1(_02979_),
    .S(_03068_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_1 _16328_ (.A(_03073_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _16329_ (.A0(net1888),
    .A1(_02981_),
    .S(_03068_),
    .X(_03074_));
 sky130_fd_sc_hd__clkbuf_1 _16330_ (.A(_03074_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _16331_ (.A0(\cur_mb_mem[126][6] ),
    .A1(_02983_),
    .S(_03068_),
    .X(_03075_));
 sky130_fd_sc_hd__clkbuf_1 _16332_ (.A(_03075_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _16333_ (.A0(net1900),
    .A1(_02985_),
    .S(_03068_),
    .X(_03076_));
 sky130_fd_sc_hd__clkbuf_1 _16334_ (.A(_03076_),
    .X(_01166_));
 sky130_fd_sc_hd__and3_1 _16335_ (.A(_02406_),
    .B(_06119_),
    .C(_03036_),
    .X(_03077_));
 sky130_fd_sc_hd__buf_4 _16336_ (.A(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__mux2_1 _16337_ (.A0(net1138),
    .A1(_02969_),
    .S(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__clkbuf_1 _16338_ (.A(_03079_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _16339_ (.A0(net1287),
    .A1(_02973_),
    .S(_03078_),
    .X(_03080_));
 sky130_fd_sc_hd__clkbuf_1 _16340_ (.A(_03080_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _16341_ (.A0(net1041),
    .A1(_02975_),
    .S(_03078_),
    .X(_03081_));
 sky130_fd_sc_hd__clkbuf_1 _16342_ (.A(_03081_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _16343_ (.A0(net1102),
    .A1(_02977_),
    .S(_03078_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_1 _16344_ (.A(_03082_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _16345_ (.A0(net970),
    .A1(_02979_),
    .S(_03078_),
    .X(_03083_));
 sky130_fd_sc_hd__clkbuf_1 _16346_ (.A(_03083_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _16347_ (.A0(net1594),
    .A1(_02981_),
    .S(_03078_),
    .X(_03084_));
 sky130_fd_sc_hd__clkbuf_1 _16348_ (.A(_03084_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _16349_ (.A0(net858),
    .A1(_02983_),
    .S(_03078_),
    .X(_03085_));
 sky130_fd_sc_hd__clkbuf_1 _16350_ (.A(_03085_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _16351_ (.A0(net876),
    .A1(_02985_),
    .S(_03078_),
    .X(_03086_));
 sky130_fd_sc_hd__clkbuf_1 _16352_ (.A(_03086_),
    .X(_01174_));
 sky130_fd_sc_hd__buf_12 _16353_ (.A(_09132_),
    .X(_03087_));
 sky130_fd_sc_hd__nand2_4 _16354_ (.A(_05935_),
    .B(_08883_),
    .Y(_03088_));
 sky130_fd_sc_hd__mux2_1 _16355_ (.A0(_03087_),
    .A1(net1285),
    .S(_03088_),
    .X(_03089_));
 sky130_fd_sc_hd__clkbuf_1 _16356_ (.A(_03089_),
    .X(_01175_));
 sky130_fd_sc_hd__clkbuf_8 _16357_ (.A(_09136_),
    .X(_03090_));
 sky130_fd_sc_hd__mux2_1 _16358_ (.A0(_03090_),
    .A1(net1864),
    .S(_03088_),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_1 _16359_ (.A(_03091_),
    .X(_01176_));
 sky130_fd_sc_hd__buf_8 _16360_ (.A(_09139_),
    .X(_03092_));
 sky130_fd_sc_hd__mux2_1 _16361_ (.A0(_03092_),
    .A1(net1549),
    .S(_03088_),
    .X(_03093_));
 sky130_fd_sc_hd__clkbuf_1 _16362_ (.A(_03093_),
    .X(_01177_));
 sky130_fd_sc_hd__clkbuf_16 _16363_ (.A(_09142_),
    .X(_03094_));
 sky130_fd_sc_hd__mux2_1 _16364_ (.A0(_03094_),
    .A1(net1686),
    .S(_03088_),
    .X(_03095_));
 sky130_fd_sc_hd__clkbuf_1 _16365_ (.A(_03095_),
    .X(_01178_));
 sky130_fd_sc_hd__buf_8 _16366_ (.A(_09145_),
    .X(_03096_));
 sky130_fd_sc_hd__mux2_1 _16367_ (.A0(_03096_),
    .A1(net1636),
    .S(_03088_),
    .X(_03097_));
 sky130_fd_sc_hd__clkbuf_1 _16368_ (.A(_03097_),
    .X(_01179_));
 sky130_fd_sc_hd__buf_8 _16369_ (.A(_09148_),
    .X(_03098_));
 sky130_fd_sc_hd__mux2_1 _16370_ (.A0(_03098_),
    .A1(net1336),
    .S(_03088_),
    .X(_03099_));
 sky130_fd_sc_hd__clkbuf_1 _16371_ (.A(_03099_),
    .X(_01180_));
 sky130_fd_sc_hd__clkbuf_8 _16372_ (.A(_09151_),
    .X(_03100_));
 sky130_fd_sc_hd__mux2_1 _16373_ (.A0(_03100_),
    .A1(net1513),
    .S(_03088_),
    .X(_03101_));
 sky130_fd_sc_hd__clkbuf_1 _16374_ (.A(_03101_),
    .X(_01181_));
 sky130_fd_sc_hd__clkbuf_8 _16375_ (.A(_09154_),
    .X(_03102_));
 sky130_fd_sc_hd__mux2_1 _16376_ (.A0(_03102_),
    .A1(net1947),
    .S(_03088_),
    .X(_03103_));
 sky130_fd_sc_hd__clkbuf_1 _16377_ (.A(_03103_),
    .X(_01182_));
 sky130_fd_sc_hd__nand2_8 _16378_ (.A(_05966_),
    .B(_02552_),
    .Y(_03104_));
 sky130_fd_sc_hd__mux2_1 _16379_ (.A0(_03087_),
    .A1(net1174),
    .S(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__clkbuf_1 _16380_ (.A(_03105_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _16381_ (.A0(_03090_),
    .A1(net1521),
    .S(_03104_),
    .X(_03106_));
 sky130_fd_sc_hd__clkbuf_1 _16382_ (.A(_03106_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _16383_ (.A0(_03092_),
    .A1(net1584),
    .S(_03104_),
    .X(_03107_));
 sky130_fd_sc_hd__clkbuf_1 _16384_ (.A(_03107_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _16385_ (.A0(_03094_),
    .A1(net1429),
    .S(_03104_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_1 _16386_ (.A(_03108_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _16387_ (.A0(_03096_),
    .A1(net733),
    .S(_03104_),
    .X(_03109_));
 sky130_fd_sc_hd__clkbuf_1 _16388_ (.A(_03109_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _16389_ (.A0(_03098_),
    .A1(net936),
    .S(_03104_),
    .X(_03110_));
 sky130_fd_sc_hd__clkbuf_1 _16390_ (.A(_03110_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _16391_ (.A0(_03100_),
    .A1(net1792),
    .S(_03104_),
    .X(_03111_));
 sky130_fd_sc_hd__clkbuf_1 _16392_ (.A(_03111_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _16393_ (.A0(_03102_),
    .A1(net1932),
    .S(_03104_),
    .X(_03112_));
 sky130_fd_sc_hd__clkbuf_1 _16394_ (.A(_03112_),
    .X(_01190_));
 sky130_fd_sc_hd__buf_12 _16395_ (.A(_08958_),
    .X(_03113_));
 sky130_fd_sc_hd__nand2_8 _16396_ (.A(_06266_),
    .B(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__mux2_1 _16397_ (.A0(_03087_),
    .A1(net607),
    .S(_03114_),
    .X(_03115_));
 sky130_fd_sc_hd__clkbuf_1 _16398_ (.A(_03115_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _16399_ (.A0(_03090_),
    .A1(net956),
    .S(_03114_),
    .X(_03116_));
 sky130_fd_sc_hd__clkbuf_1 _16400_ (.A(_03116_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _16401_ (.A0(_03092_),
    .A1(net971),
    .S(_03114_),
    .X(_03117_));
 sky130_fd_sc_hd__clkbuf_1 _16402_ (.A(_03117_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _16403_ (.A0(_03094_),
    .A1(net1022),
    .S(_03114_),
    .X(_03118_));
 sky130_fd_sc_hd__clkbuf_1 _16404_ (.A(_03118_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _16405_ (.A0(_03096_),
    .A1(net782),
    .S(_03114_),
    .X(_03119_));
 sky130_fd_sc_hd__clkbuf_1 _16406_ (.A(_03119_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _16407_ (.A0(_03098_),
    .A1(net776),
    .S(_03114_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_1 _16408_ (.A(_03120_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _16409_ (.A0(_03100_),
    .A1(net1179),
    .S(_03114_),
    .X(_03121_));
 sky130_fd_sc_hd__clkbuf_1 _16410_ (.A(_03121_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _16411_ (.A0(_03102_),
    .A1(net1707),
    .S(_03114_),
    .X(_03122_));
 sky130_fd_sc_hd__clkbuf_1 _16412_ (.A(_03122_),
    .X(_01198_));
 sky130_fd_sc_hd__nand2_8 _16413_ (.A(_06383_),
    .B(_03113_),
    .Y(_03123_));
 sky130_fd_sc_hd__mux2_1 _16414_ (.A0(_03087_),
    .A1(net1995),
    .S(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__clkbuf_1 _16415_ (.A(_03124_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _16416_ (.A0(_03090_),
    .A1(net731),
    .S(_03123_),
    .X(_03125_));
 sky130_fd_sc_hd__clkbuf_1 _16417_ (.A(_03125_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _16418_ (.A0(_03092_),
    .A1(\cur_mb_mem[131][2] ),
    .S(_03123_),
    .X(_03126_));
 sky130_fd_sc_hd__clkbuf_1 _16419_ (.A(_03126_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _16420_ (.A0(_03094_),
    .A1(net1943),
    .S(_03123_),
    .X(_03127_));
 sky130_fd_sc_hd__clkbuf_1 _16421_ (.A(_03127_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _16422_ (.A0(_03096_),
    .A1(net1001),
    .S(_03123_),
    .X(_03128_));
 sky130_fd_sc_hd__clkbuf_1 _16423_ (.A(_03128_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _16424_ (.A0(_03098_),
    .A1(net811),
    .S(_03123_),
    .X(_03129_));
 sky130_fd_sc_hd__clkbuf_1 _16425_ (.A(_03129_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _16426_ (.A0(_03100_),
    .A1(net1510),
    .S(_03123_),
    .X(_03130_));
 sky130_fd_sc_hd__clkbuf_1 _16427_ (.A(_03130_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _16428_ (.A0(_03102_),
    .A1(net1860),
    .S(_03123_),
    .X(_03131_));
 sky130_fd_sc_hd__clkbuf_1 _16429_ (.A(_03131_),
    .X(_01206_));
 sky130_fd_sc_hd__nand2_8 _16430_ (.A(net220),
    .B(_03113_),
    .Y(_03132_));
 sky130_fd_sc_hd__mux2_1 _16431_ (.A0(_03087_),
    .A1(net1086),
    .S(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__clkbuf_1 _16432_ (.A(_03133_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _16433_ (.A0(_03090_),
    .A1(net673),
    .S(_03132_),
    .X(_03134_));
 sky130_fd_sc_hd__clkbuf_1 _16434_ (.A(_03134_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _16435_ (.A0(_03092_),
    .A1(net1245),
    .S(_03132_),
    .X(_03135_));
 sky130_fd_sc_hd__clkbuf_1 _16436_ (.A(_03135_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _16437_ (.A0(_03094_),
    .A1(net1302),
    .S(_03132_),
    .X(_03136_));
 sky130_fd_sc_hd__clkbuf_1 _16438_ (.A(_03136_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _16439_ (.A0(_03096_),
    .A1(\cur_mb_mem[132][4] ),
    .S(_03132_),
    .X(_03137_));
 sky130_fd_sc_hd__clkbuf_1 _16440_ (.A(_03137_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _16441_ (.A0(_03098_),
    .A1(\cur_mb_mem[132][5] ),
    .S(_03132_),
    .X(_03138_));
 sky130_fd_sc_hd__clkbuf_1 _16442_ (.A(_03138_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _16443_ (.A0(_03100_),
    .A1(net1643),
    .S(_03132_),
    .X(_03139_));
 sky130_fd_sc_hd__clkbuf_1 _16444_ (.A(_03139_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _16445_ (.A0(_03102_),
    .A1(net1450),
    .S(_03132_),
    .X(_03140_));
 sky130_fd_sc_hd__clkbuf_1 _16446_ (.A(_03140_),
    .X(_01214_));
 sky130_fd_sc_hd__nand2_8 _16447_ (.A(_06148_),
    .B(_03113_),
    .Y(_03141_));
 sky130_fd_sc_hd__mux2_1 _16448_ (.A0(_03087_),
    .A1(net1367),
    .S(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__clkbuf_1 _16449_ (.A(_03142_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _16450_ (.A0(_03090_),
    .A1(net962),
    .S(_03141_),
    .X(_03143_));
 sky130_fd_sc_hd__clkbuf_1 _16451_ (.A(_03143_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _16452_ (.A0(_03092_),
    .A1(net724),
    .S(_03141_),
    .X(_03144_));
 sky130_fd_sc_hd__clkbuf_1 _16453_ (.A(_03144_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _16454_ (.A0(_03094_),
    .A1(net747),
    .S(_03141_),
    .X(_03145_));
 sky130_fd_sc_hd__clkbuf_1 _16455_ (.A(_03145_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _16456_ (.A0(_03096_),
    .A1(\cur_mb_mem[133][4] ),
    .S(_03141_),
    .X(_03146_));
 sky130_fd_sc_hd__clkbuf_1 _16457_ (.A(_03146_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _16458_ (.A0(_03098_),
    .A1(\cur_mb_mem[133][5] ),
    .S(_03141_),
    .X(_03147_));
 sky130_fd_sc_hd__clkbuf_1 _16459_ (.A(_03147_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _16460_ (.A0(_03100_),
    .A1(net1408),
    .S(_03141_),
    .X(_03148_));
 sky130_fd_sc_hd__clkbuf_1 _16461_ (.A(_03148_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _16462_ (.A0(_03102_),
    .A1(\cur_mb_mem[133][7] ),
    .S(_03141_),
    .X(_03149_));
 sky130_fd_sc_hd__clkbuf_1 _16463_ (.A(_03149_),
    .X(_01222_));
 sky130_fd_sc_hd__nand2_8 _16464_ (.A(_06211_),
    .B(_03113_),
    .Y(_03150_));
 sky130_fd_sc_hd__mux2_1 _16465_ (.A0(_03087_),
    .A1(\cur_mb_mem[134][0] ),
    .S(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__clkbuf_1 _16466_ (.A(_03151_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _16467_ (.A0(_03090_),
    .A1(net1441),
    .S(_03150_),
    .X(_03152_));
 sky130_fd_sc_hd__clkbuf_1 _16468_ (.A(_03152_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _16469_ (.A0(_03092_),
    .A1(net1685),
    .S(_03150_),
    .X(_03153_));
 sky130_fd_sc_hd__clkbuf_1 _16470_ (.A(_03153_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _16471_ (.A0(_03094_),
    .A1(\cur_mb_mem[134][3] ),
    .S(_03150_),
    .X(_03154_));
 sky130_fd_sc_hd__clkbuf_1 _16472_ (.A(_03154_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _16473_ (.A0(_03096_),
    .A1(net593),
    .S(_03150_),
    .X(_03155_));
 sky130_fd_sc_hd__clkbuf_1 _16474_ (.A(_03155_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _16475_ (.A0(_03098_),
    .A1(net662),
    .S(_03150_),
    .X(_03156_));
 sky130_fd_sc_hd__clkbuf_1 _16476_ (.A(_03156_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _16477_ (.A0(_03100_),
    .A1(net1609),
    .S(_03150_),
    .X(_03157_));
 sky130_fd_sc_hd__clkbuf_1 _16478_ (.A(_03157_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _16479_ (.A0(_03102_),
    .A1(\cur_mb_mem[134][7] ),
    .S(_03150_),
    .X(_03158_));
 sky130_fd_sc_hd__clkbuf_1 _16480_ (.A(_03158_),
    .X(_01230_));
 sky130_fd_sc_hd__nand2_4 _16481_ (.A(_06462_),
    .B(_03113_),
    .Y(_03159_));
 sky130_fd_sc_hd__mux2_1 _16482_ (.A0(_03087_),
    .A1(net1862),
    .S(_03159_),
    .X(_03160_));
 sky130_fd_sc_hd__clkbuf_1 _16483_ (.A(_03160_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _16484_ (.A0(_03090_),
    .A1(net788),
    .S(_03159_),
    .X(_03161_));
 sky130_fd_sc_hd__clkbuf_1 _16485_ (.A(_03161_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _16486_ (.A0(_03092_),
    .A1(net1848),
    .S(_03159_),
    .X(_03162_));
 sky130_fd_sc_hd__clkbuf_1 _16487_ (.A(_03162_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _16488_ (.A0(_03094_),
    .A1(net1692),
    .S(_03159_),
    .X(_03163_));
 sky130_fd_sc_hd__clkbuf_1 _16489_ (.A(_03163_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _16490_ (.A0(_03096_),
    .A1(net1390),
    .S(_03159_),
    .X(_03164_));
 sky130_fd_sc_hd__clkbuf_1 _16491_ (.A(_03164_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _16492_ (.A0(_03098_),
    .A1(net1365),
    .S(_03159_),
    .X(_03165_));
 sky130_fd_sc_hd__clkbuf_1 _16493_ (.A(_03165_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _16494_ (.A0(_03100_),
    .A1(\cur_mb_mem[135][6] ),
    .S(_03159_),
    .X(_03166_));
 sky130_fd_sc_hd__clkbuf_1 _16495_ (.A(_03166_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _16496_ (.A0(_03102_),
    .A1(net1815),
    .S(_03159_),
    .X(_03167_));
 sky130_fd_sc_hd__clkbuf_1 _16497_ (.A(_03167_),
    .X(_01238_));
 sky130_fd_sc_hd__nand2_8 _16498_ (.A(_06292_),
    .B(_03113_),
    .Y(_03168_));
 sky130_fd_sc_hd__mux2_1 _16499_ (.A0(_03087_),
    .A1(net562),
    .S(_03168_),
    .X(_03169_));
 sky130_fd_sc_hd__clkbuf_1 _16500_ (.A(_03169_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _16501_ (.A0(_03090_),
    .A1(net595),
    .S(_03168_),
    .X(_03170_));
 sky130_fd_sc_hd__clkbuf_1 _16502_ (.A(_03170_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _16503_ (.A0(_03092_),
    .A1(net1322),
    .S(_03168_),
    .X(_03171_));
 sky130_fd_sc_hd__clkbuf_1 _16504_ (.A(_03171_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _16505_ (.A0(_03094_),
    .A1(net664),
    .S(_03168_),
    .X(_03172_));
 sky130_fd_sc_hd__clkbuf_1 _16506_ (.A(_03172_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _16507_ (.A0(_03096_),
    .A1(net1681),
    .S(_03168_),
    .X(_03173_));
 sky130_fd_sc_hd__clkbuf_1 _16508_ (.A(_03173_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _16509_ (.A0(_03098_),
    .A1(net1583),
    .S(_03168_),
    .X(_03174_));
 sky130_fd_sc_hd__clkbuf_1 _16510_ (.A(_03174_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _16511_ (.A0(_03100_),
    .A1(net1652),
    .S(_03168_),
    .X(_03175_));
 sky130_fd_sc_hd__clkbuf_1 _16512_ (.A(_03175_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _16513_ (.A0(_03102_),
    .A1(net1508),
    .S(_03168_),
    .X(_03176_));
 sky130_fd_sc_hd__clkbuf_1 _16514_ (.A(_03176_),
    .X(_01246_));
 sky130_fd_sc_hd__nand2_8 _16515_ (.A(_05936_),
    .B(_03113_),
    .Y(_03177_));
 sky130_fd_sc_hd__mux2_1 _16516_ (.A0(_03087_),
    .A1(net568),
    .S(_03177_),
    .X(_03178_));
 sky130_fd_sc_hd__clkbuf_1 _16517_ (.A(_03178_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _16518_ (.A0(_03090_),
    .A1(net520),
    .S(_03177_),
    .X(_03179_));
 sky130_fd_sc_hd__clkbuf_1 _16519_ (.A(_03179_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _16520_ (.A0(_03092_),
    .A1(net1029),
    .S(_03177_),
    .X(_03180_));
 sky130_fd_sc_hd__clkbuf_1 _16521_ (.A(_03180_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _16522_ (.A0(_03094_),
    .A1(net596),
    .S(_03177_),
    .X(_03181_));
 sky130_fd_sc_hd__clkbuf_1 _16523_ (.A(_03181_),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _16524_ (.A0(_03096_),
    .A1(net821),
    .S(_03177_),
    .X(_03182_));
 sky130_fd_sc_hd__clkbuf_1 _16525_ (.A(_03182_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _16526_ (.A0(_03098_),
    .A1(net687),
    .S(_03177_),
    .X(_03183_));
 sky130_fd_sc_hd__clkbuf_1 _16527_ (.A(_03183_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _16528_ (.A0(_03100_),
    .A1(net1481),
    .S(_03177_),
    .X(_03184_));
 sky130_fd_sc_hd__clkbuf_1 _16529_ (.A(_03184_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _16530_ (.A0(_03102_),
    .A1(net1239),
    .S(_03177_),
    .X(_03185_));
 sky130_fd_sc_hd__clkbuf_1 _16531_ (.A(_03185_),
    .X(_01254_));
 sky130_fd_sc_hd__buf_8 _16532_ (.A(_09132_),
    .X(_03186_));
 sky130_fd_sc_hd__nand2_8 _16533_ (.A(_05934_),
    .B(_03113_),
    .Y(_03187_));
 sky130_fd_sc_hd__mux2_1 _16534_ (.A0(_03186_),
    .A1(net1289),
    .S(_03187_),
    .X(_03188_));
 sky130_fd_sc_hd__clkbuf_1 _16535_ (.A(_03188_),
    .X(_01255_));
 sky130_fd_sc_hd__clkbuf_8 _16536_ (.A(_09136_),
    .X(_03189_));
 sky130_fd_sc_hd__mux2_1 _16537_ (.A0(_03189_),
    .A1(net399),
    .S(_03187_),
    .X(_03190_));
 sky130_fd_sc_hd__clkbuf_1 _16538_ (.A(_03190_),
    .X(_01256_));
 sky130_fd_sc_hd__buf_8 _16539_ (.A(_09139_),
    .X(_03191_));
 sky130_fd_sc_hd__mux2_1 _16540_ (.A0(_03191_),
    .A1(net1354),
    .S(_03187_),
    .X(_03192_));
 sky130_fd_sc_hd__clkbuf_1 _16541_ (.A(_03192_),
    .X(_01257_));
 sky130_fd_sc_hd__buf_8 _16542_ (.A(_09142_),
    .X(_03193_));
 sky130_fd_sc_hd__mux2_1 _16543_ (.A0(_03193_),
    .A1(net1214),
    .S(_03187_),
    .X(_03194_));
 sky130_fd_sc_hd__clkbuf_1 _16544_ (.A(_03194_),
    .X(_01258_));
 sky130_fd_sc_hd__buf_8 _16545_ (.A(_09145_),
    .X(_03195_));
 sky130_fd_sc_hd__mux2_1 _16546_ (.A0(_03195_),
    .A1(net926),
    .S(_03187_),
    .X(_03196_));
 sky130_fd_sc_hd__clkbuf_1 _16547_ (.A(_03196_),
    .X(_01259_));
 sky130_fd_sc_hd__buf_8 _16548_ (.A(_09148_),
    .X(_03197_));
 sky130_fd_sc_hd__mux2_1 _16549_ (.A0(_03197_),
    .A1(net825),
    .S(_03187_),
    .X(_03198_));
 sky130_fd_sc_hd__clkbuf_1 _16550_ (.A(_03198_),
    .X(_01260_));
 sky130_fd_sc_hd__clkbuf_8 _16551_ (.A(_09151_),
    .X(_03199_));
 sky130_fd_sc_hd__mux2_1 _16552_ (.A0(_03199_),
    .A1(net1858),
    .S(_03187_),
    .X(_03200_));
 sky130_fd_sc_hd__clkbuf_1 _16553_ (.A(_03200_),
    .X(_01261_));
 sky130_fd_sc_hd__clkbuf_8 _16554_ (.A(_09154_),
    .X(_03201_));
 sky130_fd_sc_hd__mux2_1 _16555_ (.A0(_03201_),
    .A1(net1158),
    .S(_03187_),
    .X(_03202_));
 sky130_fd_sc_hd__clkbuf_1 _16556_ (.A(_03202_),
    .X(_01262_));
 sky130_fd_sc_hd__nand2_8 _16557_ (.A(_06388_),
    .B(_03113_),
    .Y(_03203_));
 sky130_fd_sc_hd__mux2_1 _16558_ (.A0(_03186_),
    .A1(net627),
    .S(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__clkbuf_1 _16559_ (.A(_03204_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _16560_ (.A0(_03189_),
    .A1(net1257),
    .S(_03203_),
    .X(_03205_));
 sky130_fd_sc_hd__clkbuf_1 _16561_ (.A(_03205_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _16562_ (.A0(_03191_),
    .A1(net1241),
    .S(_03203_),
    .X(_03206_));
 sky130_fd_sc_hd__clkbuf_1 _16563_ (.A(_03206_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _16564_ (.A0(_03193_),
    .A1(net608),
    .S(_03203_),
    .X(_03207_));
 sky130_fd_sc_hd__clkbuf_1 _16565_ (.A(_03207_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _16566_ (.A0(_03195_),
    .A1(net830),
    .S(_03203_),
    .X(_03208_));
 sky130_fd_sc_hd__clkbuf_1 _16567_ (.A(_03208_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _16568_ (.A0(_03197_),
    .A1(net1129),
    .S(_03203_),
    .X(_03209_));
 sky130_fd_sc_hd__clkbuf_1 _16569_ (.A(_03209_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _16570_ (.A0(_03199_),
    .A1(net1353),
    .S(_03203_),
    .X(_03210_));
 sky130_fd_sc_hd__clkbuf_1 _16571_ (.A(_03210_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _16572_ (.A0(_03201_),
    .A1(net1299),
    .S(_03203_),
    .X(_03211_));
 sky130_fd_sc_hd__clkbuf_1 _16573_ (.A(_03211_),
    .X(_01270_));
 sky130_fd_sc_hd__buf_12 _16574_ (.A(_08958_),
    .X(_03212_));
 sky130_fd_sc_hd__nand2_8 _16575_ (.A(_06423_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__mux2_1 _16576_ (.A0(_03186_),
    .A1(net1605),
    .S(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__clkbuf_1 _16577_ (.A(_03214_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _16578_ (.A0(_03189_),
    .A1(net709),
    .S(_03213_),
    .X(_03215_));
 sky130_fd_sc_hd__clkbuf_1 _16579_ (.A(_03215_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _16580_ (.A0(_03191_),
    .A1(net1097),
    .S(_03213_),
    .X(_03216_));
 sky130_fd_sc_hd__clkbuf_1 _16581_ (.A(_03216_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _16582_ (.A0(_03193_),
    .A1(net1757),
    .S(_03213_),
    .X(_03217_));
 sky130_fd_sc_hd__clkbuf_1 _16583_ (.A(_03217_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _16584_ (.A0(_03195_),
    .A1(net1461),
    .S(_03213_),
    .X(_03218_));
 sky130_fd_sc_hd__clkbuf_1 _16585_ (.A(_03218_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _16586_ (.A0(_03197_),
    .A1(net1306),
    .S(_03213_),
    .X(_03219_));
 sky130_fd_sc_hd__clkbuf_1 _16587_ (.A(_03219_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _16588_ (.A0(_03199_),
    .A1(net1471),
    .S(_03213_),
    .X(_03220_));
 sky130_fd_sc_hd__clkbuf_1 _16589_ (.A(_03220_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _16590_ (.A0(_03201_),
    .A1(net1507),
    .S(_03213_),
    .X(_03221_));
 sky130_fd_sc_hd__clkbuf_1 _16591_ (.A(_03221_),
    .X(_01278_));
 sky130_fd_sc_hd__nand2_8 _16592_ (.A(_06250_),
    .B(_03212_),
    .Y(_03222_));
 sky130_fd_sc_hd__mux2_1 _16593_ (.A0(_03186_),
    .A1(net1333),
    .S(_03222_),
    .X(_03223_));
 sky130_fd_sc_hd__clkbuf_1 _16594_ (.A(_03223_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _16595_ (.A0(_03189_),
    .A1(net1372),
    .S(_03222_),
    .X(_03224_));
 sky130_fd_sc_hd__clkbuf_1 _16596_ (.A(_03224_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _16597_ (.A0(_03191_),
    .A1(net1434),
    .S(_03222_),
    .X(_03225_));
 sky130_fd_sc_hd__clkbuf_1 _16598_ (.A(_03225_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _16599_ (.A0(_03193_),
    .A1(net1135),
    .S(_03222_),
    .X(_03226_));
 sky130_fd_sc_hd__clkbuf_1 _16600_ (.A(_03226_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _16601_ (.A0(_03195_),
    .A1(net927),
    .S(_03222_),
    .X(_03227_));
 sky130_fd_sc_hd__clkbuf_1 _16602_ (.A(_03227_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _16603_ (.A0(_03197_),
    .A1(net1059),
    .S(_03222_),
    .X(_03228_));
 sky130_fd_sc_hd__clkbuf_1 _16604_ (.A(_03228_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _16605_ (.A0(_03199_),
    .A1(net1242),
    .S(_03222_),
    .X(_03229_));
 sky130_fd_sc_hd__clkbuf_1 _16606_ (.A(_03229_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _16607_ (.A0(_03201_),
    .A1(net1268),
    .S(_03222_),
    .X(_03230_));
 sky130_fd_sc_hd__clkbuf_1 _16608_ (.A(_03230_),
    .X(_01286_));
 sky130_fd_sc_hd__nand2_8 _16609_ (.A(_06487_),
    .B(_03212_),
    .Y(_03231_));
 sky130_fd_sc_hd__mux2_1 _16610_ (.A0(_03186_),
    .A1(net1165),
    .S(_03231_),
    .X(_03232_));
 sky130_fd_sc_hd__clkbuf_1 _16611_ (.A(_03232_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _16612_ (.A0(_03189_),
    .A1(net1324),
    .S(_03231_),
    .X(_03233_));
 sky130_fd_sc_hd__clkbuf_1 _16613_ (.A(_03233_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _16614_ (.A0(_03191_),
    .A1(net1342),
    .S(_03231_),
    .X(_03234_));
 sky130_fd_sc_hd__clkbuf_1 _16615_ (.A(_03234_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _16616_ (.A0(_03193_),
    .A1(net1406),
    .S(_03231_),
    .X(_03235_));
 sky130_fd_sc_hd__clkbuf_1 _16617_ (.A(_03235_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _16618_ (.A0(_03195_),
    .A1(net632),
    .S(_03231_),
    .X(_03236_));
 sky130_fd_sc_hd__clkbuf_1 _16619_ (.A(_03236_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _16620_ (.A0(_03197_),
    .A1(net726),
    .S(_03231_),
    .X(_03237_));
 sky130_fd_sc_hd__clkbuf_1 _16621_ (.A(_03237_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _16622_ (.A0(_03199_),
    .A1(net1814),
    .S(_03231_),
    .X(_03238_));
 sky130_fd_sc_hd__clkbuf_1 _16623_ (.A(_03238_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _16624_ (.A0(_03201_),
    .A1(net1816),
    .S(_03231_),
    .X(_03239_));
 sky130_fd_sc_hd__clkbuf_1 _16625_ (.A(_03239_),
    .X(_01294_));
 sky130_fd_sc_hd__nand2_8 _16626_ (.A(_06305_),
    .B(_03212_),
    .Y(_03240_));
 sky130_fd_sc_hd__mux2_1 _16627_ (.A0(_03186_),
    .A1(net1598),
    .S(_03240_),
    .X(_03241_));
 sky130_fd_sc_hd__clkbuf_1 _16628_ (.A(_03241_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _16629_ (.A0(_03189_),
    .A1(net1323),
    .S(_03240_),
    .X(_03242_));
 sky130_fd_sc_hd__clkbuf_1 _16630_ (.A(_03242_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _16631_ (.A0(_03191_),
    .A1(net1624),
    .S(_03240_),
    .X(_03243_));
 sky130_fd_sc_hd__clkbuf_1 _16632_ (.A(_03243_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _16633_ (.A0(_03193_),
    .A1(net1668),
    .S(_03240_),
    .X(_03244_));
 sky130_fd_sc_hd__clkbuf_1 _16634_ (.A(_03244_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _16635_ (.A0(_03195_),
    .A1(net1021),
    .S(_03240_),
    .X(_03245_));
 sky130_fd_sc_hd__clkbuf_1 _16636_ (.A(_03245_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _16637_ (.A0(_03197_),
    .A1(net1420),
    .S(_03240_),
    .X(_03246_));
 sky130_fd_sc_hd__clkbuf_1 _16638_ (.A(_03246_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _16639_ (.A0(_03199_),
    .A1(net1222),
    .S(_03240_),
    .X(_03247_));
 sky130_fd_sc_hd__clkbuf_1 _16640_ (.A(_03247_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _16641_ (.A0(_03201_),
    .A1(net1527),
    .S(_03240_),
    .X(_03248_));
 sky130_fd_sc_hd__clkbuf_1 _16642_ (.A(_03248_),
    .X(_01302_));
 sky130_fd_sc_hd__buf_4 _16643_ (.A(_05980_),
    .X(_03249_));
 sky130_fd_sc_hd__nand2_8 _16644_ (.A(_03249_),
    .B(_08883_),
    .Y(_03250_));
 sky130_fd_sc_hd__mux2_1 _16645_ (.A0(_03186_),
    .A1(net1619),
    .S(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__clkbuf_1 _16646_ (.A(_03251_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _16647_ (.A0(_03189_),
    .A1(net965),
    .S(_03250_),
    .X(_03252_));
 sky130_fd_sc_hd__clkbuf_1 _16648_ (.A(_03252_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _16649_ (.A0(_03191_),
    .A1(net1637),
    .S(_03250_),
    .X(_03253_));
 sky130_fd_sc_hd__clkbuf_1 _16650_ (.A(_03253_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _16651_ (.A0(_03193_),
    .A1(net1642),
    .S(_03250_),
    .X(_03254_));
 sky130_fd_sc_hd__clkbuf_1 _16652_ (.A(_03254_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _16653_ (.A0(_03195_),
    .A1(net666),
    .S(_03250_),
    .X(_03255_));
 sky130_fd_sc_hd__clkbuf_1 _16654_ (.A(_03255_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _16655_ (.A0(_03197_),
    .A1(net765),
    .S(_03250_),
    .X(_03256_));
 sky130_fd_sc_hd__clkbuf_1 _16656_ (.A(_03256_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _16657_ (.A0(_03199_),
    .A1(net1156),
    .S(_03250_),
    .X(_03257_));
 sky130_fd_sc_hd__clkbuf_1 _16658_ (.A(_03257_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _16659_ (.A0(_03201_),
    .A1(net1081),
    .S(_03250_),
    .X(_03258_));
 sky130_fd_sc_hd__clkbuf_1 _16660_ (.A(_03258_),
    .X(_01310_));
 sky130_fd_sc_hd__nand2_8 _16661_ (.A(_06252_),
    .B(_03212_),
    .Y(_03259_));
 sky130_fd_sc_hd__mux2_1 _16662_ (.A0(_03186_),
    .A1(net781),
    .S(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__clkbuf_1 _16663_ (.A(_03260_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _16664_ (.A0(_03189_),
    .A1(net1430),
    .S(_03259_),
    .X(_03261_));
 sky130_fd_sc_hd__clkbuf_1 _16665_ (.A(_03261_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _16666_ (.A0(_03191_),
    .A1(net1200),
    .S(_03259_),
    .X(_03262_));
 sky130_fd_sc_hd__clkbuf_1 _16667_ (.A(_03262_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _16668_ (.A0(_03193_),
    .A1(net570),
    .S(_03259_),
    .X(_03263_));
 sky130_fd_sc_hd__clkbuf_1 _16669_ (.A(_03263_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _16670_ (.A0(_03195_),
    .A1(net745),
    .S(_03259_),
    .X(_03264_));
 sky130_fd_sc_hd__clkbuf_1 _16671_ (.A(_03264_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _16672_ (.A0(_03197_),
    .A1(net1110),
    .S(_03259_),
    .X(_03265_));
 sky130_fd_sc_hd__clkbuf_1 _16673_ (.A(_03265_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _16674_ (.A0(_03199_),
    .A1(net1217),
    .S(_03259_),
    .X(_03266_));
 sky130_fd_sc_hd__clkbuf_1 _16675_ (.A(_03266_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _16676_ (.A0(_03201_),
    .A1(net1272),
    .S(_03259_),
    .X(_03267_));
 sky130_fd_sc_hd__clkbuf_1 _16677_ (.A(_03267_),
    .X(_01318_));
 sky130_fd_sc_hd__nand2_8 _16678_ (.A(_06381_),
    .B(_03212_),
    .Y(_03268_));
 sky130_fd_sc_hd__mux2_1 _16679_ (.A0(_03186_),
    .A1(net798),
    .S(_03268_),
    .X(_03269_));
 sky130_fd_sc_hd__clkbuf_1 _16680_ (.A(_03269_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _16681_ (.A0(_03189_),
    .A1(net451),
    .S(_03268_),
    .X(_03270_));
 sky130_fd_sc_hd__clkbuf_1 _16682_ (.A(_03270_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _16683_ (.A0(_03191_),
    .A1(net989),
    .S(_03268_),
    .X(_03271_));
 sky130_fd_sc_hd__clkbuf_1 _16684_ (.A(_03271_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _16685_ (.A0(_03193_),
    .A1(net1093),
    .S(_03268_),
    .X(_03272_));
 sky130_fd_sc_hd__clkbuf_1 _16686_ (.A(_03272_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _16687_ (.A0(_03195_),
    .A1(net1183),
    .S(_03268_),
    .X(_03273_));
 sky130_fd_sc_hd__clkbuf_1 _16688_ (.A(_03273_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _16689_ (.A0(_03197_),
    .A1(net1485),
    .S(_03268_),
    .X(_03274_));
 sky130_fd_sc_hd__clkbuf_1 _16690_ (.A(_03274_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _16691_ (.A0(_03199_),
    .A1(net1447),
    .S(_03268_),
    .X(_03275_));
 sky130_fd_sc_hd__clkbuf_1 _16692_ (.A(_03275_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _16693_ (.A0(_03201_),
    .A1(net1867),
    .S(_03268_),
    .X(_03276_));
 sky130_fd_sc_hd__clkbuf_1 _16694_ (.A(_03276_),
    .X(_01326_));
 sky130_fd_sc_hd__buf_8 _16695_ (.A(_08530_),
    .X(_03277_));
 sky130_fd_sc_hd__and3_1 _16696_ (.A(_02266_),
    .B(_03249_),
    .C(_03036_),
    .X(_03278_));
 sky130_fd_sc_hd__buf_8 _16697_ (.A(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__mux2_1 _16698_ (.A0(net535),
    .A1(_03277_),
    .S(_03279_),
    .X(_03280_));
 sky130_fd_sc_hd__clkbuf_1 _16699_ (.A(_03280_),
    .X(_01327_));
 sky130_fd_sc_hd__buf_4 _16700_ (.A(_08535_),
    .X(_03281_));
 sky130_fd_sc_hd__mux2_1 _16701_ (.A0(net350),
    .A1(_03281_),
    .S(_03279_),
    .X(_03282_));
 sky130_fd_sc_hd__clkbuf_1 _16702_ (.A(_03282_),
    .X(_01328_));
 sky130_fd_sc_hd__clkbuf_8 _16703_ (.A(_08538_),
    .X(_03283_));
 sky130_fd_sc_hd__mux2_1 _16704_ (.A0(net1026),
    .A1(_03283_),
    .S(_03279_),
    .X(_03284_));
 sky130_fd_sc_hd__clkbuf_1 _16705_ (.A(_03284_),
    .X(_01329_));
 sky130_fd_sc_hd__clkbuf_8 _16706_ (.A(_08541_),
    .X(_03285_));
 sky130_fd_sc_hd__mux2_1 _16707_ (.A0(net680),
    .A1(_03285_),
    .S(_03279_),
    .X(_03286_));
 sky130_fd_sc_hd__clkbuf_1 _16708_ (.A(_03286_),
    .X(_01330_));
 sky130_fd_sc_hd__clkbuf_4 _16709_ (.A(_08544_),
    .X(_03287_));
 sky130_fd_sc_hd__mux2_1 _16710_ (.A0(net1491),
    .A1(_03287_),
    .S(_03279_),
    .X(_03288_));
 sky130_fd_sc_hd__clkbuf_1 _16711_ (.A(_03288_),
    .X(_01331_));
 sky130_fd_sc_hd__buf_4 _16712_ (.A(_08547_),
    .X(_03289_));
 sky130_fd_sc_hd__mux2_1 _16713_ (.A0(net1618),
    .A1(_03289_),
    .S(_03279_),
    .X(_03290_));
 sky130_fd_sc_hd__clkbuf_1 _16714_ (.A(_03290_),
    .X(_01332_));
 sky130_fd_sc_hd__clkbuf_8 _16715_ (.A(_08550_),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_1 _16716_ (.A0(net445),
    .A1(_03291_),
    .S(_03279_),
    .X(_03292_));
 sky130_fd_sc_hd__clkbuf_1 _16717_ (.A(_03292_),
    .X(_01333_));
 sky130_fd_sc_hd__buf_4 _16718_ (.A(_08553_),
    .X(_03293_));
 sky130_fd_sc_hd__mux2_1 _16719_ (.A0(net759),
    .A1(_03293_),
    .S(_03279_),
    .X(_03294_));
 sky130_fd_sc_hd__clkbuf_1 _16720_ (.A(_03294_),
    .X(_01334_));
 sky130_fd_sc_hd__nand3_4 _16721_ (.A(_06223_),
    .B(_03249_),
    .C(_08901_),
    .Y(_03295_));
 sky130_fd_sc_hd__mux2_1 _16722_ (.A0(_03186_),
    .A1(net1855),
    .S(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__clkbuf_1 _16723_ (.A(_03296_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _16724_ (.A0(_03189_),
    .A1(net646),
    .S(_03295_),
    .X(_03297_));
 sky130_fd_sc_hd__clkbuf_1 _16725_ (.A(_03297_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _16726_ (.A0(_03191_),
    .A1(net1807),
    .S(_03295_),
    .X(_03298_));
 sky130_fd_sc_hd__clkbuf_1 _16727_ (.A(_03298_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _16728_ (.A0(_03193_),
    .A1(net1826),
    .S(_03295_),
    .X(_03299_));
 sky130_fd_sc_hd__clkbuf_1 _16729_ (.A(_03299_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _16730_ (.A0(_03195_),
    .A1(net843),
    .S(_03295_),
    .X(_03300_));
 sky130_fd_sc_hd__clkbuf_1 _16731_ (.A(_03300_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _16732_ (.A0(_03197_),
    .A1(net581),
    .S(_03295_),
    .X(_03301_));
 sky130_fd_sc_hd__clkbuf_1 _16733_ (.A(_03301_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _16734_ (.A0(_03199_),
    .A1(net1301),
    .S(_03295_),
    .X(_03302_));
 sky130_fd_sc_hd__clkbuf_1 _16735_ (.A(_03302_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _16736_ (.A0(_03201_),
    .A1(net1219),
    .S(_03295_),
    .X(_03303_));
 sky130_fd_sc_hd__clkbuf_1 _16737_ (.A(_03303_),
    .X(_01342_));
 sky130_fd_sc_hd__and3_1 _16738_ (.A(_03249_),
    .B(_02286_),
    .C(_03036_),
    .X(_03304_));
 sky130_fd_sc_hd__buf_4 _16739_ (.A(_03304_),
    .X(_03305_));
 sky130_fd_sc_hd__mux2_1 _16740_ (.A0(net1115),
    .A1(_03277_),
    .S(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__clkbuf_1 _16741_ (.A(_03306_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _16742_ (.A0(net633),
    .A1(_03281_),
    .S(_03305_),
    .X(_03307_));
 sky130_fd_sc_hd__clkbuf_1 _16743_ (.A(_03307_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _16744_ (.A0(net1410),
    .A1(_03283_),
    .S(_03305_),
    .X(_03308_));
 sky130_fd_sc_hd__clkbuf_1 _16745_ (.A(_03308_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _16746_ (.A0(net510),
    .A1(_03285_),
    .S(_03305_),
    .X(_03309_));
 sky130_fd_sc_hd__clkbuf_1 _16747_ (.A(_03309_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _16748_ (.A0(net552),
    .A1(_03287_),
    .S(_03305_),
    .X(_03310_));
 sky130_fd_sc_hd__clkbuf_1 _16749_ (.A(_03310_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _16750_ (.A0(net502),
    .A1(_03289_),
    .S(_03305_),
    .X(_03311_));
 sky130_fd_sc_hd__clkbuf_1 _16751_ (.A(_03311_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _16752_ (.A0(\cur_mb_mem[149][6] ),
    .A1(_03291_),
    .S(_03305_),
    .X(_03312_));
 sky130_fd_sc_hd__clkbuf_1 _16753_ (.A(_03312_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _16754_ (.A0(net816),
    .A1(_03293_),
    .S(_03305_),
    .X(_03313_));
 sky130_fd_sc_hd__clkbuf_1 _16755_ (.A(_03313_),
    .X(_01350_));
 sky130_fd_sc_hd__and3_1 _16756_ (.A(_02297_),
    .B(_03249_),
    .C(_03036_),
    .X(_03314_));
 sky130_fd_sc_hd__clkbuf_8 _16757_ (.A(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__mux2_1 _16758_ (.A0(net584),
    .A1(_03277_),
    .S(_03315_),
    .X(_03316_));
 sky130_fd_sc_hd__clkbuf_1 _16759_ (.A(_03316_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _16760_ (.A0(net853),
    .A1(_03281_),
    .S(_03315_),
    .X(_03317_));
 sky130_fd_sc_hd__clkbuf_1 _16761_ (.A(_03317_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _16762_ (.A0(net1123),
    .A1(_03283_),
    .S(_03315_),
    .X(_03318_));
 sky130_fd_sc_hd__clkbuf_1 _16763_ (.A(_03318_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _16764_ (.A0(net1327),
    .A1(_03285_),
    .S(_03315_),
    .X(_03319_));
 sky130_fd_sc_hd__clkbuf_1 _16765_ (.A(_03319_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _16766_ (.A0(net966),
    .A1(_03287_),
    .S(_03315_),
    .X(_03320_));
 sky130_fd_sc_hd__clkbuf_1 _16767_ (.A(_03320_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _16768_ (.A0(net1262),
    .A1(_03289_),
    .S(_03315_),
    .X(_03321_));
 sky130_fd_sc_hd__clkbuf_1 _16769_ (.A(_03321_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _16770_ (.A0(net1610),
    .A1(_03291_),
    .S(_03315_),
    .X(_03322_));
 sky130_fd_sc_hd__clkbuf_1 _16771_ (.A(_03322_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _16772_ (.A0(net893),
    .A1(_03293_),
    .S(_03315_),
    .X(_03323_));
 sky130_fd_sc_hd__clkbuf_1 _16773_ (.A(_03323_),
    .X(_01358_));
 sky130_fd_sc_hd__and3_1 _16774_ (.A(_03249_),
    .B(_08839_),
    .C(_03036_),
    .X(_03324_));
 sky130_fd_sc_hd__clkbuf_8 _16775_ (.A(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__mux2_1 _16776_ (.A0(net1620),
    .A1(_03277_),
    .S(_03325_),
    .X(_03326_));
 sky130_fd_sc_hd__clkbuf_1 _16777_ (.A(_03326_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _16778_ (.A0(net981),
    .A1(_03281_),
    .S(_03325_),
    .X(_03327_));
 sky130_fd_sc_hd__clkbuf_1 _16779_ (.A(_03327_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _16780_ (.A0(net1851),
    .A1(_03283_),
    .S(_03325_),
    .X(_03328_));
 sky130_fd_sc_hd__clkbuf_1 _16781_ (.A(_03328_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _16782_ (.A0(net1615),
    .A1(_03285_),
    .S(_03325_),
    .X(_03329_));
 sky130_fd_sc_hd__clkbuf_1 _16783_ (.A(_03329_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _16784_ (.A0(net1253),
    .A1(_03287_),
    .S(_03325_),
    .X(_03330_));
 sky130_fd_sc_hd__clkbuf_1 _16785_ (.A(_03330_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _16786_ (.A0(net1495),
    .A1(_03289_),
    .S(_03325_),
    .X(_03331_));
 sky130_fd_sc_hd__clkbuf_1 _16787_ (.A(_03331_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _16788_ (.A0(net1885),
    .A1(_03291_),
    .S(_03325_),
    .X(_03332_));
 sky130_fd_sc_hd__clkbuf_1 _16789_ (.A(_03332_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _16790_ (.A0(net1256),
    .A1(_03293_),
    .S(_03325_),
    .X(_03333_));
 sky130_fd_sc_hd__clkbuf_1 _16791_ (.A(_03333_),
    .X(_01366_));
 sky130_fd_sc_hd__clkbuf_16 _16792_ (.A(_09132_),
    .X(_03334_));
 sky130_fd_sc_hd__nand2_8 _16793_ (.A(_06394_),
    .B(_03212_),
    .Y(_03335_));
 sky130_fd_sc_hd__mux2_1 _16794_ (.A0(_03334_),
    .A1(net1341),
    .S(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__clkbuf_1 _16795_ (.A(_03336_),
    .X(_01367_));
 sky130_fd_sc_hd__buf_6 _16796_ (.A(_09136_),
    .X(_03337_));
 sky130_fd_sc_hd__mux2_1 _16797_ (.A0(_03337_),
    .A1(net1356),
    .S(_03335_),
    .X(_03338_));
 sky130_fd_sc_hd__clkbuf_1 _16798_ (.A(_03338_),
    .X(_01368_));
 sky130_fd_sc_hd__buf_8 _16799_ (.A(_09139_),
    .X(_03339_));
 sky130_fd_sc_hd__mux2_1 _16800_ (.A0(_03339_),
    .A1(net1100),
    .S(_03335_),
    .X(_03340_));
 sky130_fd_sc_hd__clkbuf_1 _16801_ (.A(_03340_),
    .X(_01369_));
 sky130_fd_sc_hd__buf_8 _16802_ (.A(_09142_),
    .X(_03341_));
 sky130_fd_sc_hd__mux2_1 _16803_ (.A0(_03341_),
    .A1(net1586),
    .S(_03335_),
    .X(_03342_));
 sky130_fd_sc_hd__clkbuf_1 _16804_ (.A(_03342_),
    .X(_01370_));
 sky130_fd_sc_hd__clkbuf_16 _16805_ (.A(_09145_),
    .X(_03343_));
 sky130_fd_sc_hd__mux2_1 _16806_ (.A0(_03343_),
    .A1(net1313),
    .S(_03335_),
    .X(_03344_));
 sky130_fd_sc_hd__clkbuf_1 _16807_ (.A(_03344_),
    .X(_01371_));
 sky130_fd_sc_hd__buf_12 _16808_ (.A(_09148_),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_1 _16809_ (.A0(_03345_),
    .A1(net1276),
    .S(_03335_),
    .X(_03346_));
 sky130_fd_sc_hd__clkbuf_1 _16810_ (.A(_03346_),
    .X(_01372_));
 sky130_fd_sc_hd__clkbuf_8 _16811_ (.A(_09151_),
    .X(_03347_));
 sky130_fd_sc_hd__mux2_1 _16812_ (.A0(_03347_),
    .A1(net1109),
    .S(_03335_),
    .X(_03348_));
 sky130_fd_sc_hd__clkbuf_1 _16813_ (.A(_03348_),
    .X(_01373_));
 sky130_fd_sc_hd__clkbuf_8 _16814_ (.A(_09154_),
    .X(_03349_));
 sky130_fd_sc_hd__mux2_1 _16815_ (.A0(_03349_),
    .A1(net1706),
    .S(_03335_),
    .X(_03350_));
 sky130_fd_sc_hd__clkbuf_1 _16816_ (.A(_03350_),
    .X(_01374_));
 sky130_fd_sc_hd__and3_1 _16817_ (.A(_08978_),
    .B(_03249_),
    .C(_03036_),
    .X(_03351_));
 sky130_fd_sc_hd__buf_4 _16818_ (.A(_03351_),
    .X(_03352_));
 sky130_fd_sc_hd__mux2_1 _16819_ (.A0(net450),
    .A1(_03277_),
    .S(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__clkbuf_1 _16820_ (.A(_03353_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _16821_ (.A0(net1778),
    .A1(_03281_),
    .S(_03352_),
    .X(_03354_));
 sky130_fd_sc_hd__clkbuf_1 _16822_ (.A(_03354_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _16823_ (.A0(net313),
    .A1(_03283_),
    .S(_03352_),
    .X(_03355_));
 sky130_fd_sc_hd__clkbuf_1 _16824_ (.A(_03355_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _16825_ (.A0(net441),
    .A1(_03285_),
    .S(_03352_),
    .X(_03356_));
 sky130_fd_sc_hd__clkbuf_1 _16826_ (.A(_03356_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _16827_ (.A0(net1601),
    .A1(_03287_),
    .S(_03352_),
    .X(_03357_));
 sky130_fd_sc_hd__clkbuf_1 _16828_ (.A(_03357_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _16829_ (.A0(net1772),
    .A1(_03289_),
    .S(_03352_),
    .X(_03358_));
 sky130_fd_sc_hd__clkbuf_1 _16830_ (.A(_03358_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _16831_ (.A0(\cur_mb_mem[153][6] ),
    .A1(_03291_),
    .S(_03352_),
    .X(_03359_));
 sky130_fd_sc_hd__clkbuf_1 _16832_ (.A(_03359_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _16833_ (.A0(\cur_mb_mem[153][7] ),
    .A1(_03293_),
    .S(_03352_),
    .X(_03360_));
 sky130_fd_sc_hd__clkbuf_1 _16834_ (.A(_03360_),
    .X(_01382_));
 sky130_fd_sc_hd__clkbuf_4 _16835_ (.A(_08900_),
    .X(_03361_));
 sky130_fd_sc_hd__and3_1 _16836_ (.A(_02353_),
    .B(_03249_),
    .C(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__buf_4 _16837_ (.A(_03362_),
    .X(_03363_));
 sky130_fd_sc_hd__mux2_1 _16838_ (.A0(net1494),
    .A1(_03277_),
    .S(_03363_),
    .X(_03364_));
 sky130_fd_sc_hd__clkbuf_1 _16839_ (.A(_03364_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _16840_ (.A0(net1781),
    .A1(_03281_),
    .S(_03363_),
    .X(_03365_));
 sky130_fd_sc_hd__clkbuf_1 _16841_ (.A(_03365_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _16842_ (.A0(net372),
    .A1(_03283_),
    .S(_03363_),
    .X(_03366_));
 sky130_fd_sc_hd__clkbuf_1 _16843_ (.A(_03366_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _16844_ (.A0(net458),
    .A1(_03285_),
    .S(_03363_),
    .X(_03367_));
 sky130_fd_sc_hd__clkbuf_1 _16845_ (.A(_03367_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _16846_ (.A0(net1451),
    .A1(_03287_),
    .S(_03363_),
    .X(_03368_));
 sky130_fd_sc_hd__clkbuf_1 _16847_ (.A(_03368_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _16848_ (.A0(net1409),
    .A1(_03289_),
    .S(_03363_),
    .X(_03369_));
 sky130_fd_sc_hd__clkbuf_1 _16849_ (.A(_03369_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _16850_ (.A0(net972),
    .A1(_03291_),
    .S(_03363_),
    .X(_03370_));
 sky130_fd_sc_hd__clkbuf_1 _16851_ (.A(_03370_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _16852_ (.A0(net931),
    .A1(_03293_),
    .S(_03363_),
    .X(_03371_));
 sky130_fd_sc_hd__clkbuf_1 _16853_ (.A(_03371_),
    .X(_01390_));
 sky130_fd_sc_hd__and3_1 _16854_ (.A(_02526_),
    .B(_03249_),
    .C(_03361_),
    .X(_03372_));
 sky130_fd_sc_hd__buf_4 _16855_ (.A(_03372_),
    .X(_03373_));
 sky130_fd_sc_hd__mux2_1 _16856_ (.A0(net1820),
    .A1(_03277_),
    .S(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__clkbuf_1 _16857_ (.A(_03374_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _16858_ (.A0(net339),
    .A1(_03281_),
    .S(_03373_),
    .X(_03375_));
 sky130_fd_sc_hd__clkbuf_1 _16859_ (.A(_03375_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _16860_ (.A0(net1237),
    .A1(_03283_),
    .S(_03373_),
    .X(_03376_));
 sky130_fd_sc_hd__clkbuf_1 _16861_ (.A(_03376_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _16862_ (.A0(net1743),
    .A1(_03285_),
    .S(_03373_),
    .X(_03377_));
 sky130_fd_sc_hd__clkbuf_1 _16863_ (.A(_03377_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _16864_ (.A0(net1189),
    .A1(_03287_),
    .S(_03373_),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_1 _16865_ (.A(_03378_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _16866_ (.A0(net763),
    .A1(_03289_),
    .S(_03373_),
    .X(_03379_));
 sky130_fd_sc_hd__clkbuf_1 _16867_ (.A(_03379_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _16868_ (.A0(\cur_mb_mem[155][6] ),
    .A1(_03291_),
    .S(_03373_),
    .X(_03380_));
 sky130_fd_sc_hd__clkbuf_1 _16869_ (.A(_03380_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _16870_ (.A0(net1942),
    .A1(_03293_),
    .S(_03373_),
    .X(_03381_));
 sky130_fd_sc_hd__clkbuf_1 _16871_ (.A(_03381_),
    .X(_01398_));
 sky130_fd_sc_hd__and3_1 _16872_ (.A(_02374_),
    .B(_05980_),
    .C(_03361_),
    .X(_03382_));
 sky130_fd_sc_hd__buf_4 _16873_ (.A(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__mux2_1 _16874_ (.A0(net1879),
    .A1(_03277_),
    .S(_03383_),
    .X(_03384_));
 sky130_fd_sc_hd__clkbuf_1 _16875_ (.A(_03384_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _16876_ (.A0(net919),
    .A1(_03281_),
    .S(_03383_),
    .X(_03385_));
 sky130_fd_sc_hd__clkbuf_1 _16877_ (.A(_03385_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _16878_ (.A0(net1710),
    .A1(_03283_),
    .S(_03383_),
    .X(_03386_));
 sky130_fd_sc_hd__clkbuf_1 _16879_ (.A(_03386_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _16880_ (.A0(net1722),
    .A1(_03285_),
    .S(_03383_),
    .X(_03387_));
 sky130_fd_sc_hd__clkbuf_1 _16881_ (.A(_03387_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _16882_ (.A0(net921),
    .A1(_03287_),
    .S(_03383_),
    .X(_03388_));
 sky130_fd_sc_hd__clkbuf_1 _16883_ (.A(_03388_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _16884_ (.A0(net852),
    .A1(_03289_),
    .S(_03383_),
    .X(_03389_));
 sky130_fd_sc_hd__clkbuf_1 _16885_ (.A(_03389_),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _16886_ (.A0(net1213),
    .A1(_03291_),
    .S(_03383_),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_1 _16887_ (.A(_03390_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _16888_ (.A0(net803),
    .A1(_03293_),
    .S(_03383_),
    .X(_03391_));
 sky130_fd_sc_hd__clkbuf_1 _16889_ (.A(_03391_),
    .X(_01406_));
 sky130_fd_sc_hd__and3_1 _16890_ (.A(_09025_),
    .B(_05980_),
    .C(_03361_),
    .X(_03392_));
 sky130_fd_sc_hd__buf_6 _16891_ (.A(_03392_),
    .X(_03393_));
 sky130_fd_sc_hd__mux2_1 _16892_ (.A0(net1504),
    .A1(_03277_),
    .S(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__clkbuf_1 _16893_ (.A(_03394_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _16894_ (.A0(net424),
    .A1(_03281_),
    .S(_03393_),
    .X(_03395_));
 sky130_fd_sc_hd__clkbuf_1 _16895_ (.A(_03395_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _16896_ (.A0(net1641),
    .A1(_03283_),
    .S(_03393_),
    .X(_03396_));
 sky130_fd_sc_hd__clkbuf_1 _16897_ (.A(_03396_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _16898_ (.A0(net819),
    .A1(_03285_),
    .S(_03393_),
    .X(_03397_));
 sky130_fd_sc_hd__clkbuf_1 _16899_ (.A(_03397_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _16900_ (.A0(net1645),
    .A1(_03287_),
    .S(_03393_),
    .X(_03398_));
 sky130_fd_sc_hd__clkbuf_1 _16901_ (.A(_03398_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _16902_ (.A0(net1563),
    .A1(_03289_),
    .S(_03393_),
    .X(_03399_));
 sky130_fd_sc_hd__clkbuf_1 _16903_ (.A(_03399_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _16904_ (.A0(net1033),
    .A1(_03291_),
    .S(_03393_),
    .X(_03400_));
 sky130_fd_sc_hd__clkbuf_1 _16905_ (.A(_03400_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _16906_ (.A0(net1014),
    .A1(_03293_),
    .S(_03393_),
    .X(_03401_));
 sky130_fd_sc_hd__clkbuf_1 _16907_ (.A(_03401_),
    .X(_01414_));
 sky130_fd_sc_hd__and3_1 _16908_ (.A(_03249_),
    .B(_09036_),
    .C(_03361_),
    .X(_03402_));
 sky130_fd_sc_hd__buf_4 _16909_ (.A(_03402_),
    .X(_03403_));
 sky130_fd_sc_hd__mux2_1 _16910_ (.A0(net428),
    .A1(_03277_),
    .S(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_1 _16911_ (.A(_03404_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _16912_ (.A0(net1013),
    .A1(_03281_),
    .S(_03403_),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_1 _16913_ (.A(_03405_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _16914_ (.A0(net1401),
    .A1(_03283_),
    .S(_03403_),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_1 _16915_ (.A(_03406_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _16916_ (.A0(net401),
    .A1(_03285_),
    .S(_03403_),
    .X(_03407_));
 sky130_fd_sc_hd__clkbuf_1 _16917_ (.A(_03407_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _16918_ (.A0(net1416),
    .A1(_03287_),
    .S(_03403_),
    .X(_03408_));
 sky130_fd_sc_hd__clkbuf_1 _16919_ (.A(_03408_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _16920_ (.A0(net1520),
    .A1(_03289_),
    .S(_03403_),
    .X(_03409_));
 sky130_fd_sc_hd__clkbuf_1 _16921_ (.A(_03409_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _16922_ (.A0(\cur_mb_mem[158][6] ),
    .A1(_03291_),
    .S(_03403_),
    .X(_03410_));
 sky130_fd_sc_hd__clkbuf_1 _16923_ (.A(_03410_),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _16924_ (.A0(net1878),
    .A1(_03293_),
    .S(_03403_),
    .X(_03411_));
 sky130_fd_sc_hd__clkbuf_1 _16925_ (.A(_03411_),
    .X(_01422_));
 sky130_fd_sc_hd__buf_12 _16926_ (.A(_08530_),
    .X(_03412_));
 sky130_fd_sc_hd__and3_1 _16927_ (.A(_02406_),
    .B(_05980_),
    .C(_03361_),
    .X(_03413_));
 sky130_fd_sc_hd__buf_6 _16928_ (.A(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__mux2_1 _16929_ (.A0(net1067),
    .A1(_03412_),
    .S(_03414_),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_1 _16930_ (.A(_03415_),
    .X(_01423_));
 sky130_fd_sc_hd__clkbuf_16 _16931_ (.A(_08535_),
    .X(_03416_));
 sky130_fd_sc_hd__mux2_1 _16932_ (.A0(net1695),
    .A1(_03416_),
    .S(_03414_),
    .X(_03417_));
 sky130_fd_sc_hd__clkbuf_1 _16933_ (.A(_03417_),
    .X(_01424_));
 sky130_fd_sc_hd__buf_12 _16934_ (.A(_08538_),
    .X(_03418_));
 sky130_fd_sc_hd__mux2_1 _16935_ (.A0(net1230),
    .A1(_03418_),
    .S(_03414_),
    .X(_03419_));
 sky130_fd_sc_hd__clkbuf_1 _16936_ (.A(_03419_),
    .X(_01425_));
 sky130_fd_sc_hd__buf_12 _16937_ (.A(_08541_),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_1 _16938_ (.A0(net1467),
    .A1(_03420_),
    .S(_03414_),
    .X(_03421_));
 sky130_fd_sc_hd__clkbuf_1 _16939_ (.A(_03421_),
    .X(_01426_));
 sky130_fd_sc_hd__buf_8 _16940_ (.A(_08544_),
    .X(_03422_));
 sky130_fd_sc_hd__mux2_1 _16941_ (.A0(net942),
    .A1(_03422_),
    .S(_03414_),
    .X(_03423_));
 sky130_fd_sc_hd__clkbuf_1 _16942_ (.A(_03423_),
    .X(_01427_));
 sky130_fd_sc_hd__buf_8 _16943_ (.A(_08547_),
    .X(_03424_));
 sky130_fd_sc_hd__mux2_1 _16944_ (.A0(net1665),
    .A1(_03424_),
    .S(_03414_),
    .X(_03425_));
 sky130_fd_sc_hd__clkbuf_1 _16945_ (.A(_03425_),
    .X(_01428_));
 sky130_fd_sc_hd__clkbuf_16 _16946_ (.A(_08550_),
    .X(_03426_));
 sky130_fd_sc_hd__mux2_1 _16947_ (.A0(net717),
    .A1(_03426_),
    .S(_03414_),
    .X(_03427_));
 sky130_fd_sc_hd__clkbuf_1 _16948_ (.A(_03427_),
    .X(_01429_));
 sky130_fd_sc_hd__buf_6 _16949_ (.A(_08553_),
    .X(_03428_));
 sky130_fd_sc_hd__mux2_1 _16950_ (.A0(net1137),
    .A1(_03428_),
    .S(_03414_),
    .X(_03429_));
 sky130_fd_sc_hd__clkbuf_1 _16951_ (.A(_03429_),
    .X(_01430_));
 sky130_fd_sc_hd__buf_4 _16952_ (.A(_05956_),
    .X(_03430_));
 sky130_fd_sc_hd__nand2_8 _16953_ (.A(_03430_),
    .B(_08882_),
    .Y(_03431_));
 sky130_fd_sc_hd__mux2_1 _16954_ (.A0(_03334_),
    .A1(net889),
    .S(_03431_),
    .X(_03432_));
 sky130_fd_sc_hd__clkbuf_1 _16955_ (.A(_03432_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _16956_ (.A0(_03337_),
    .A1(net1056),
    .S(_03431_),
    .X(_03433_));
 sky130_fd_sc_hd__clkbuf_1 _16957_ (.A(_03433_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _16958_ (.A0(_03339_),
    .A1(net1403),
    .S(_03431_),
    .X(_03434_));
 sky130_fd_sc_hd__clkbuf_1 _16959_ (.A(_03434_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _16960_ (.A0(_03341_),
    .A1(net1018),
    .S(_03431_),
    .X(_03435_));
 sky130_fd_sc_hd__clkbuf_1 _16961_ (.A(_03435_),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _16962_ (.A0(_03343_),
    .A1(net637),
    .S(_03431_),
    .X(_03436_));
 sky130_fd_sc_hd__clkbuf_1 _16963_ (.A(_03436_),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _16964_ (.A0(_03345_),
    .A1(net547),
    .S(_03431_),
    .X(_03437_));
 sky130_fd_sc_hd__clkbuf_1 _16965_ (.A(_03437_),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _16966_ (.A0(_03347_),
    .A1(net1448),
    .S(_03431_),
    .X(_03438_));
 sky130_fd_sc_hd__clkbuf_1 _16967_ (.A(_03438_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _16968_ (.A0(_03349_),
    .A1(net555),
    .S(_03431_),
    .X(_03439_));
 sky130_fd_sc_hd__clkbuf_1 _16969_ (.A(_03439_),
    .X(_01438_));
 sky130_fd_sc_hd__nand2_8 _16970_ (.A(_06334_),
    .B(_03212_),
    .Y(_03440_));
 sky130_fd_sc_hd__mux2_1 _16971_ (.A0(_03334_),
    .A1(net1411),
    .S(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__clkbuf_1 _16972_ (.A(_03441_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _16973_ (.A0(_03337_),
    .A1(net1087),
    .S(_03440_),
    .X(_03442_));
 sky130_fd_sc_hd__clkbuf_1 _16974_ (.A(_03442_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _16975_ (.A0(_03339_),
    .A1(net1582),
    .S(_03440_),
    .X(_03443_));
 sky130_fd_sc_hd__clkbuf_1 _16976_ (.A(_03443_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _16977_ (.A0(_03341_),
    .A1(net1140),
    .S(_03440_),
    .X(_03444_));
 sky130_fd_sc_hd__clkbuf_1 _16978_ (.A(_03444_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _16979_ (.A0(_03343_),
    .A1(net866),
    .S(_03440_),
    .X(_03445_));
 sky130_fd_sc_hd__clkbuf_1 _16980_ (.A(_03445_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _16981_ (.A0(_03345_),
    .A1(net1019),
    .S(_03440_),
    .X(_03446_));
 sky130_fd_sc_hd__clkbuf_1 _16982_ (.A(_03446_),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _16983_ (.A0(_03347_),
    .A1(net1455),
    .S(_03440_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_1 _16984_ (.A(_03447_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _16985_ (.A0(_03349_),
    .A1(net1194),
    .S(_03440_),
    .X(_03448_));
 sky130_fd_sc_hd__clkbuf_1 _16986_ (.A(_03448_),
    .X(_01446_));
 sky130_fd_sc_hd__nand2_8 _16987_ (.A(_06284_),
    .B(_03212_),
    .Y(_03449_));
 sky130_fd_sc_hd__mux2_1 _16988_ (.A0(_03334_),
    .A1(net820),
    .S(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__clkbuf_1 _16989_ (.A(_03450_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _16990_ (.A0(_03337_),
    .A1(net621),
    .S(_03449_),
    .X(_03451_));
 sky130_fd_sc_hd__clkbuf_1 _16991_ (.A(_03451_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _16992_ (.A0(_03339_),
    .A1(net1201),
    .S(_03449_),
    .X(_03452_));
 sky130_fd_sc_hd__clkbuf_1 _16993_ (.A(_03452_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _16994_ (.A0(_03341_),
    .A1(net834),
    .S(_03449_),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_1 _16995_ (.A(_03453_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _16996_ (.A0(_03343_),
    .A1(net1474),
    .S(_03449_),
    .X(_03454_));
 sky130_fd_sc_hd__clkbuf_1 _16997_ (.A(_03454_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _16998_ (.A0(_03345_),
    .A1(net1375),
    .S(_03449_),
    .X(_03455_));
 sky130_fd_sc_hd__clkbuf_1 _16999_ (.A(_03455_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _17000_ (.A0(_03347_),
    .A1(net1112),
    .S(_03449_),
    .X(_03456_));
 sky130_fd_sc_hd__clkbuf_1 _17001_ (.A(_03456_),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _17002_ (.A0(_03349_),
    .A1(net1204),
    .S(_03449_),
    .X(_03457_));
 sky130_fd_sc_hd__clkbuf_1 _17003_ (.A(_03457_),
    .X(_01454_));
 sky130_fd_sc_hd__and3_1 _17004_ (.A(_02266_),
    .B(_03430_),
    .C(_03361_),
    .X(_03458_));
 sky130_fd_sc_hd__buf_6 _17005_ (.A(_03458_),
    .X(_03459_));
 sky130_fd_sc_hd__mux2_1 _17006_ (.A0(net484),
    .A1(_03412_),
    .S(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__clkbuf_1 _17007_ (.A(_03460_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _17008_ (.A0(net363),
    .A1(_03416_),
    .S(_03459_),
    .X(_03461_));
 sky130_fd_sc_hd__clkbuf_1 _17009_ (.A(_03461_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _17010_ (.A0(net571),
    .A1(_03418_),
    .S(_03459_),
    .X(_03462_));
 sky130_fd_sc_hd__clkbuf_1 _17011_ (.A(_03462_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _17012_ (.A0(net690),
    .A1(_03420_),
    .S(_03459_),
    .X(_03463_));
 sky130_fd_sc_hd__clkbuf_1 _17013_ (.A(_03463_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _17014_ (.A0(net550),
    .A1(_03422_),
    .S(_03459_),
    .X(_03464_));
 sky130_fd_sc_hd__clkbuf_1 _17015_ (.A(_03464_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _17016_ (.A0(net472),
    .A1(_03424_),
    .S(_03459_),
    .X(_03465_));
 sky130_fd_sc_hd__clkbuf_1 _17017_ (.A(_03465_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _17018_ (.A0(net964),
    .A1(_03426_),
    .S(_03459_),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_1 _17019_ (.A(_03466_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _17020_ (.A0(net1069),
    .A1(_03428_),
    .S(_03459_),
    .X(_03467_));
 sky130_fd_sc_hd__clkbuf_1 _17021_ (.A(_03467_),
    .X(_01462_));
 sky130_fd_sc_hd__nand2_8 _17022_ (.A(_06195_),
    .B(_03212_),
    .Y(_03468_));
 sky130_fd_sc_hd__mux2_1 _17023_ (.A0(_03334_),
    .A1(net1533),
    .S(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_1 _17024_ (.A(_03469_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _17025_ (.A0(_03337_),
    .A1(net1613),
    .S(_03468_),
    .X(_03470_));
 sky130_fd_sc_hd__clkbuf_1 _17026_ (.A(_03470_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _17027_ (.A0(_03339_),
    .A1(net1452),
    .S(_03468_),
    .X(_03471_));
 sky130_fd_sc_hd__clkbuf_1 _17028_ (.A(_03471_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _17029_ (.A0(_03341_),
    .A1(net1498),
    .S(_03468_),
    .X(_03472_));
 sky130_fd_sc_hd__clkbuf_1 _17030_ (.A(_03472_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _17031_ (.A0(_03343_),
    .A1(net1173),
    .S(_03468_),
    .X(_03473_));
 sky130_fd_sc_hd__clkbuf_1 _17032_ (.A(_03473_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _17033_ (.A0(_03345_),
    .A1(net1159),
    .S(_03468_),
    .X(_03474_));
 sky130_fd_sc_hd__clkbuf_1 _17034_ (.A(_03474_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _17035_ (.A0(_03347_),
    .A1(net1238),
    .S(_03468_),
    .X(_03475_));
 sky130_fd_sc_hd__clkbuf_1 _17036_ (.A(_03475_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _17037_ (.A0(_03349_),
    .A1(net1057),
    .S(_03468_),
    .X(_03476_));
 sky130_fd_sc_hd__clkbuf_1 _17038_ (.A(_03476_),
    .X(_01470_));
 sky130_fd_sc_hd__and3_1 _17039_ (.A(_03430_),
    .B(_02286_),
    .C(_03361_),
    .X(_03477_));
 sky130_fd_sc_hd__buf_8 _17040_ (.A(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__mux2_1 _17041_ (.A0(net417),
    .A1(_03412_),
    .S(_03478_),
    .X(_03479_));
 sky130_fd_sc_hd__clkbuf_1 _17042_ (.A(_03479_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _17043_ (.A0(net352),
    .A1(_03416_),
    .S(_03478_),
    .X(_03480_));
 sky130_fd_sc_hd__clkbuf_1 _17044_ (.A(_03480_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _17045_ (.A0(net325),
    .A1(_03418_),
    .S(_03478_),
    .X(_03481_));
 sky130_fd_sc_hd__clkbuf_1 _17046_ (.A(_03481_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _17047_ (.A0(net758),
    .A1(_03420_),
    .S(_03478_),
    .X(_03482_));
 sky130_fd_sc_hd__clkbuf_1 _17048_ (.A(_03482_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _17049_ (.A0(net660),
    .A1(_03422_),
    .S(_03478_),
    .X(_03483_));
 sky130_fd_sc_hd__clkbuf_1 _17050_ (.A(_03483_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _17051_ (.A0(net409),
    .A1(_03424_),
    .S(_03478_),
    .X(_03484_));
 sky130_fd_sc_hd__clkbuf_1 _17052_ (.A(_03484_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _17053_ (.A0(net995),
    .A1(_03426_),
    .S(_03478_),
    .X(_03485_));
 sky130_fd_sc_hd__clkbuf_1 _17054_ (.A(_03485_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _17055_ (.A0(net1380),
    .A1(_03428_),
    .S(_03478_),
    .X(_03486_));
 sky130_fd_sc_hd__clkbuf_1 _17056_ (.A(_03486_),
    .X(_01478_));
 sky130_fd_sc_hd__and3_1 _17057_ (.A(_02297_),
    .B(_03430_),
    .C(_03361_),
    .X(_03487_));
 sky130_fd_sc_hd__buf_6 _17058_ (.A(_03487_),
    .X(_03488_));
 sky130_fd_sc_hd__mux2_1 _17059_ (.A0(net1075),
    .A1(_03412_),
    .S(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__clkbuf_1 _17060_ (.A(_03489_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _17061_ (.A0(net780),
    .A1(_03416_),
    .S(_03488_),
    .X(_03490_));
 sky130_fd_sc_hd__clkbuf_1 _17062_ (.A(_03490_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _17063_ (.A0(net986),
    .A1(_03418_),
    .S(_03488_),
    .X(_03491_));
 sky130_fd_sc_hd__clkbuf_1 _17064_ (.A(_03491_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _17065_ (.A0(net1361),
    .A1(_03420_),
    .S(_03488_),
    .X(_03492_));
 sky130_fd_sc_hd__clkbuf_1 _17066_ (.A(_03492_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _17067_ (.A0(net1125),
    .A1(_03422_),
    .S(_03488_),
    .X(_03493_));
 sky130_fd_sc_hd__clkbuf_1 _17068_ (.A(_03493_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _17069_ (.A0(net1180),
    .A1(_03424_),
    .S(_03488_),
    .X(_03494_));
 sky130_fd_sc_hd__clkbuf_1 _17070_ (.A(_03494_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _17071_ (.A0(net1167),
    .A1(_03426_),
    .S(_03488_),
    .X(_03495_));
 sky130_fd_sc_hd__clkbuf_1 _17072_ (.A(_03495_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _17073_ (.A0(net880),
    .A1(_03428_),
    .S(_03488_),
    .X(_03496_));
 sky130_fd_sc_hd__clkbuf_1 _17074_ (.A(_03496_),
    .X(_01486_));
 sky130_fd_sc_hd__and3_1 _17075_ (.A(_03430_),
    .B(_08839_),
    .C(_03361_),
    .X(_03497_));
 sky130_fd_sc_hd__buf_4 _17076_ (.A(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__mux2_1 _17077_ (.A0(net556),
    .A1(_03412_),
    .S(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__clkbuf_1 _17078_ (.A(_03499_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _17079_ (.A0(net485),
    .A1(_03416_),
    .S(_03498_),
    .X(_03500_));
 sky130_fd_sc_hd__clkbuf_1 _17080_ (.A(_03500_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _17081_ (.A0(net509),
    .A1(_03418_),
    .S(_03498_),
    .X(_03501_));
 sky130_fd_sc_hd__clkbuf_1 _17082_ (.A(_03501_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _17083_ (.A0(net421),
    .A1(_03420_),
    .S(_03498_),
    .X(_03502_));
 sky130_fd_sc_hd__clkbuf_1 _17084_ (.A(_03502_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _17085_ (.A0(net1186),
    .A1(_03422_),
    .S(_03498_),
    .X(_03503_));
 sky130_fd_sc_hd__clkbuf_1 _17086_ (.A(_03503_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _17087_ (.A0(net1344),
    .A1(_03424_),
    .S(_03498_),
    .X(_03504_));
 sky130_fd_sc_hd__clkbuf_1 _17088_ (.A(_03504_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _17089_ (.A0(net940),
    .A1(_03426_),
    .S(_03498_),
    .X(_03505_));
 sky130_fd_sc_hd__clkbuf_1 _17090_ (.A(_03505_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _17091_ (.A0(net1037),
    .A1(_03428_),
    .S(_03498_),
    .X(_03506_));
 sky130_fd_sc_hd__clkbuf_1 _17092_ (.A(_03506_),
    .X(_01494_));
 sky130_fd_sc_hd__nand3_4 _17093_ (.A(_05896_),
    .B(_03430_),
    .C(_08901_),
    .Y(_03507_));
 sky130_fd_sc_hd__mux2_1 _17094_ (.A0(_03334_),
    .A1(net592),
    .S(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__clkbuf_1 _17095_ (.A(_03508_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _17096_ (.A0(_03337_),
    .A1(net1025),
    .S(_03507_),
    .X(_03509_));
 sky130_fd_sc_hd__clkbuf_1 _17097_ (.A(_03509_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _17098_ (.A0(_03339_),
    .A1(net767),
    .S(_03507_),
    .X(_03510_));
 sky130_fd_sc_hd__clkbuf_1 _17099_ (.A(_03510_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _17100_ (.A0(_03341_),
    .A1(net1338),
    .S(_03507_),
    .X(_03511_));
 sky130_fd_sc_hd__clkbuf_1 _17101_ (.A(_03511_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _17102_ (.A0(_03343_),
    .A1(net760),
    .S(_03507_),
    .X(_03512_));
 sky130_fd_sc_hd__clkbuf_1 _17103_ (.A(_03512_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _17104_ (.A0(_03345_),
    .A1(net1902),
    .S(_03507_),
    .X(_03513_));
 sky130_fd_sc_hd__clkbuf_1 _17105_ (.A(_03513_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _17106_ (.A0(_03347_),
    .A1(net1445),
    .S(_03507_),
    .X(_03514_));
 sky130_fd_sc_hd__clkbuf_1 _17107_ (.A(_03514_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _17108_ (.A0(_03349_),
    .A1(net1465),
    .S(_03507_),
    .X(_03515_));
 sky130_fd_sc_hd__clkbuf_1 _17109_ (.A(_03515_),
    .X(_01502_));
 sky130_fd_sc_hd__buf_2 _17110_ (.A(_08900_),
    .X(_03516_));
 sky130_fd_sc_hd__and3_1 _17111_ (.A(_08978_),
    .B(_03430_),
    .C(_03516_),
    .X(_03517_));
 sky130_fd_sc_hd__buf_6 _17112_ (.A(_03517_),
    .X(_03518_));
 sky130_fd_sc_hd__mux2_1 _17113_ (.A0(net980),
    .A1(_03412_),
    .S(_03518_),
    .X(_03519_));
 sky130_fd_sc_hd__clkbuf_1 _17114_ (.A(_03519_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _17115_ (.A0(net573),
    .A1(_03416_),
    .S(_03518_),
    .X(_03520_));
 sky130_fd_sc_hd__clkbuf_1 _17116_ (.A(_03520_),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _17117_ (.A0(net448),
    .A1(_03418_),
    .S(_03518_),
    .X(_03521_));
 sky130_fd_sc_hd__clkbuf_1 _17118_ (.A(_03521_),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _17119_ (.A0(net619),
    .A1(_03420_),
    .S(_03518_),
    .X(_03522_));
 sky130_fd_sc_hd__clkbuf_1 _17120_ (.A(_03522_),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _17121_ (.A0(net503),
    .A1(_03422_),
    .S(_03518_),
    .X(_03523_));
 sky130_fd_sc_hd__clkbuf_1 _17122_ (.A(_03523_),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _17123_ (.A0(net382),
    .A1(_03424_),
    .S(_03518_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_1 _17124_ (.A(_03524_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _17125_ (.A0(net863),
    .A1(_03426_),
    .S(_03518_),
    .X(_03525_));
 sky130_fd_sc_hd__clkbuf_1 _17126_ (.A(_03525_),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _17127_ (.A0(net974),
    .A1(_03428_),
    .S(_03518_),
    .X(_03526_));
 sky130_fd_sc_hd__clkbuf_1 _17128_ (.A(_03526_),
    .X(_01510_));
 sky130_fd_sc_hd__and3_1 _17129_ (.A(_02353_),
    .B(_03430_),
    .C(_03516_),
    .X(_03527_));
 sky130_fd_sc_hd__buf_6 _17130_ (.A(_03527_),
    .X(_03528_));
 sky130_fd_sc_hd__mux2_1 _17131_ (.A0(net469),
    .A1(_03412_),
    .S(_03528_),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_1 _17132_ (.A(_03529_),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _17133_ (.A0(net774),
    .A1(_03416_),
    .S(_03528_),
    .X(_03530_));
 sky130_fd_sc_hd__clkbuf_1 _17134_ (.A(_03530_),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _17135_ (.A0(net447),
    .A1(_03418_),
    .S(_03528_),
    .X(_03531_));
 sky130_fd_sc_hd__clkbuf_1 _17136_ (.A(_03531_),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _17137_ (.A0(net321),
    .A1(_03420_),
    .S(_03528_),
    .X(_03532_));
 sky130_fd_sc_hd__clkbuf_1 _17138_ (.A(_03532_),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_1 _17139_ (.A0(net665),
    .A1(_03422_),
    .S(_03528_),
    .X(_03533_));
 sky130_fd_sc_hd__clkbuf_1 _17140_ (.A(_03533_),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _17141_ (.A0(net415),
    .A1(_03424_),
    .S(_03528_),
    .X(_03534_));
 sky130_fd_sc_hd__clkbuf_1 _17142_ (.A(_03534_),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _17143_ (.A0(net1017),
    .A1(_03426_),
    .S(_03528_),
    .X(_03535_));
 sky130_fd_sc_hd__clkbuf_1 _17144_ (.A(_03535_),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _17145_ (.A0(net314),
    .A1(_03428_),
    .S(_03528_),
    .X(_03536_));
 sky130_fd_sc_hd__clkbuf_1 _17146_ (.A(_03536_),
    .X(_01518_));
 sky130_fd_sc_hd__and3_1 _17147_ (.A(_02526_),
    .B(_03430_),
    .C(_03516_),
    .X(_03537_));
 sky130_fd_sc_hd__buf_6 _17148_ (.A(_03537_),
    .X(_03538_));
 sky130_fd_sc_hd__mux2_1 _17149_ (.A0(net383),
    .A1(_03412_),
    .S(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__clkbuf_1 _17150_ (.A(_03539_),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _17151_ (.A0(net603),
    .A1(_03416_),
    .S(_03538_),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_1 _17152_ (.A(_03540_),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _17153_ (.A0(net406),
    .A1(_03418_),
    .S(_03538_),
    .X(_03541_));
 sky130_fd_sc_hd__clkbuf_1 _17154_ (.A(_03541_),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _17155_ (.A0(net460),
    .A1(_03420_),
    .S(_03538_),
    .X(_03542_));
 sky130_fd_sc_hd__clkbuf_1 _17156_ (.A(_03542_),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _17157_ (.A0(net335),
    .A1(_03422_),
    .S(_03538_),
    .X(_03543_));
 sky130_fd_sc_hd__clkbuf_1 _17158_ (.A(_03543_),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _17159_ (.A0(net508),
    .A1(_03424_),
    .S(_03538_),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_1 _17160_ (.A(_03544_),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _17161_ (.A0(net710),
    .A1(_03426_),
    .S(_03538_),
    .X(_03545_));
 sky130_fd_sc_hd__clkbuf_1 _17162_ (.A(_03545_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _17163_ (.A0(net468),
    .A1(_03428_),
    .S(_03538_),
    .X(_03546_));
 sky130_fd_sc_hd__clkbuf_1 _17164_ (.A(_03546_),
    .X(_01526_));
 sky130_fd_sc_hd__and3_1 _17165_ (.A(_02374_),
    .B(_03430_),
    .C(_03516_),
    .X(_03547_));
 sky130_fd_sc_hd__buf_8 _17166_ (.A(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__mux2_1 _17167_ (.A0(net537),
    .A1(_03412_),
    .S(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__clkbuf_1 _17168_ (.A(_03549_),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _17169_ (.A0(net394),
    .A1(_03416_),
    .S(_03548_),
    .X(_03550_));
 sky130_fd_sc_hd__clkbuf_1 _17170_ (.A(_03550_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _17171_ (.A0(net695),
    .A1(_03418_),
    .S(_03548_),
    .X(_03551_));
 sky130_fd_sc_hd__clkbuf_1 _17172_ (.A(_03551_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _17173_ (.A0(net342),
    .A1(_03420_),
    .S(_03548_),
    .X(_03552_));
 sky130_fd_sc_hd__clkbuf_1 _17174_ (.A(_03552_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _17175_ (.A0(net443),
    .A1(_03422_),
    .S(_03548_),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_1 _17176_ (.A(_03553_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _17177_ (.A0(net505),
    .A1(_03424_),
    .S(_03548_),
    .X(_03554_));
 sky130_fd_sc_hd__clkbuf_1 _17178_ (.A(_03554_),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _17179_ (.A0(net1185),
    .A1(_03426_),
    .S(_03548_),
    .X(_03555_));
 sky130_fd_sc_hd__clkbuf_1 _17180_ (.A(_03555_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _17181_ (.A0(net899),
    .A1(_03428_),
    .S(_03548_),
    .X(_03556_));
 sky130_fd_sc_hd__clkbuf_1 _17182_ (.A(_03556_),
    .X(_01534_));
 sky130_fd_sc_hd__and3_1 _17183_ (.A(_09025_),
    .B(_05956_),
    .C(_03516_),
    .X(_03557_));
 sky130_fd_sc_hd__buf_4 _17184_ (.A(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__mux2_1 _17185_ (.A0(net403),
    .A1(_03412_),
    .S(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__clkbuf_1 _17186_ (.A(_03559_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _17187_ (.A0(net500),
    .A1(_03416_),
    .S(_03558_),
    .X(_03560_));
 sky130_fd_sc_hd__clkbuf_1 _17188_ (.A(_03560_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _17189_ (.A0(net477),
    .A1(_03418_),
    .S(_03558_),
    .X(_03561_));
 sky130_fd_sc_hd__clkbuf_1 _17190_ (.A(_03561_),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _17191_ (.A0(net525),
    .A1(_03420_),
    .S(_03558_),
    .X(_03562_));
 sky130_fd_sc_hd__clkbuf_1 _17192_ (.A(_03562_),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _17193_ (.A0(net391),
    .A1(_03422_),
    .S(_03558_),
    .X(_03563_));
 sky130_fd_sc_hd__clkbuf_1 _17194_ (.A(_03563_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _17195_ (.A0(net371),
    .A1(_03424_),
    .S(_03558_),
    .X(_03564_));
 sky130_fd_sc_hd__clkbuf_1 _17196_ (.A(_03564_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _17197_ (.A0(net1062),
    .A1(_03426_),
    .S(_03558_),
    .X(_03565_));
 sky130_fd_sc_hd__clkbuf_1 _17198_ (.A(_03565_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _17199_ (.A0(net1094),
    .A1(_03428_),
    .S(_03558_),
    .X(_03566_));
 sky130_fd_sc_hd__clkbuf_1 _17200_ (.A(_03566_),
    .X(_01542_));
 sky130_fd_sc_hd__buf_8 _17201_ (.A(_08530_),
    .X(_03567_));
 sky130_fd_sc_hd__and3_1 _17202_ (.A(_09036_),
    .B(_05956_),
    .C(_03516_),
    .X(_03568_));
 sky130_fd_sc_hd__clkbuf_8 _17203_ (.A(_03568_),
    .X(_03569_));
 sky130_fd_sc_hd__mux2_1 _17204_ (.A0(net1131),
    .A1(_03567_),
    .S(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__clkbuf_1 _17205_ (.A(_03570_),
    .X(_01543_));
 sky130_fd_sc_hd__buf_6 _17206_ (.A(_08535_),
    .X(_03571_));
 sky130_fd_sc_hd__mux2_1 _17207_ (.A0(net361),
    .A1(_03571_),
    .S(_03569_),
    .X(_03572_));
 sky130_fd_sc_hd__clkbuf_1 _17208_ (.A(_03572_),
    .X(_01544_));
 sky130_fd_sc_hd__buf_8 _17209_ (.A(_08538_),
    .X(_03573_));
 sky130_fd_sc_hd__mux2_1 _17210_ (.A0(net355),
    .A1(_03573_),
    .S(_03569_),
    .X(_03574_));
 sky130_fd_sc_hd__clkbuf_1 _17211_ (.A(_03574_),
    .X(_01545_));
 sky130_fd_sc_hd__buf_8 _17212_ (.A(_08541_),
    .X(_03575_));
 sky130_fd_sc_hd__mux2_1 _17213_ (.A0(net671),
    .A1(_03575_),
    .S(_03569_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_1 _17214_ (.A(_03576_),
    .X(_01546_));
 sky130_fd_sc_hd__buf_8 _17215_ (.A(_08544_),
    .X(_03577_));
 sky130_fd_sc_hd__mux2_1 _17216_ (.A0(net436),
    .A1(_03577_),
    .S(_03569_),
    .X(_03578_));
 sky130_fd_sc_hd__clkbuf_1 _17217_ (.A(_03578_),
    .X(_01547_));
 sky130_fd_sc_hd__buf_8 _17218_ (.A(_08547_),
    .X(_03579_));
 sky130_fd_sc_hd__mux2_1 _17219_ (.A0(net324),
    .A1(_03579_),
    .S(_03569_),
    .X(_03580_));
 sky130_fd_sc_hd__clkbuf_1 _17220_ (.A(_03580_),
    .X(_01548_));
 sky130_fd_sc_hd__clkbuf_8 _17221_ (.A(_08550_),
    .X(_03581_));
 sky130_fd_sc_hd__mux2_1 _17222_ (.A0(net845),
    .A1(_03581_),
    .S(_03569_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_1 _17223_ (.A(_03582_),
    .X(_01549_));
 sky130_fd_sc_hd__buf_4 _17224_ (.A(_08553_),
    .X(_03583_));
 sky130_fd_sc_hd__mux2_1 _17225_ (.A0(net829),
    .A1(_03583_),
    .S(_03569_),
    .X(_03584_));
 sky130_fd_sc_hd__clkbuf_1 _17226_ (.A(_03584_),
    .X(_01550_));
 sky130_fd_sc_hd__and3_1 _17227_ (.A(_02406_),
    .B(_05956_),
    .C(_03516_),
    .X(_03585_));
 sky130_fd_sc_hd__clkbuf_8 _17228_ (.A(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__mux2_1 _17229_ (.A0(net1235),
    .A1(_03567_),
    .S(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__clkbuf_1 _17230_ (.A(_03587_),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _17231_ (.A0(net539),
    .A1(_03571_),
    .S(_03586_),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_1 _17232_ (.A(_03588_),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _17233_ (.A0(net998),
    .A1(_03573_),
    .S(_03586_),
    .X(_03589_));
 sky130_fd_sc_hd__clkbuf_1 _17234_ (.A(_03589_),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _17235_ (.A0(net1319),
    .A1(_03575_),
    .S(_03586_),
    .X(_03590_));
 sky130_fd_sc_hd__clkbuf_1 _17236_ (.A(_03590_),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _17237_ (.A0(net770),
    .A1(_03577_),
    .S(_03586_),
    .X(_03591_));
 sky130_fd_sc_hd__clkbuf_1 _17238_ (.A(_03591_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _17239_ (.A0(net380),
    .A1(_03579_),
    .S(_03586_),
    .X(_03592_));
 sky130_fd_sc_hd__clkbuf_1 _17240_ (.A(_03592_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _17241_ (.A0(net842),
    .A1(_03581_),
    .S(_03586_),
    .X(_03593_));
 sky130_fd_sc_hd__clkbuf_1 _17242_ (.A(_03593_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _17243_ (.A0(net1133),
    .A1(_03583_),
    .S(_03586_),
    .X(_03594_));
 sky130_fd_sc_hd__clkbuf_1 _17244_ (.A(_03594_),
    .X(_01558_));
 sky130_fd_sc_hd__buf_4 _17245_ (.A(_06037_),
    .X(_03595_));
 sky130_fd_sc_hd__nand2_8 _17246_ (.A(_03595_),
    .B(_08882_),
    .Y(_03596_));
 sky130_fd_sc_hd__mux2_1 _17247_ (.A0(_03334_),
    .A1(net1489),
    .S(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__clkbuf_1 _17248_ (.A(_03597_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _17249_ (.A0(_03337_),
    .A1(net846),
    .S(_03596_),
    .X(_03598_));
 sky130_fd_sc_hd__clkbuf_1 _17250_ (.A(_03598_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _17251_ (.A0(_03339_),
    .A1(net1236),
    .S(_03596_),
    .X(_03599_));
 sky130_fd_sc_hd__clkbuf_1 _17252_ (.A(_03599_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _17253_ (.A0(_03341_),
    .A1(net1351),
    .S(_03596_),
    .X(_03600_));
 sky130_fd_sc_hd__clkbuf_1 _17254_ (.A(_03600_),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _17255_ (.A0(_03343_),
    .A1(net1148),
    .S(_03596_),
    .X(_03601_));
 sky130_fd_sc_hd__clkbuf_1 _17256_ (.A(_03601_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _17257_ (.A0(_03345_),
    .A1(net544),
    .S(_03596_),
    .X(_03602_));
 sky130_fd_sc_hd__clkbuf_1 _17258_ (.A(_03602_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _17259_ (.A0(_03347_),
    .A1(net1715),
    .S(_03596_),
    .X(_03603_));
 sky130_fd_sc_hd__clkbuf_1 _17260_ (.A(_03603_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _17261_ (.A0(_03349_),
    .A1(net1177),
    .S(_03596_),
    .X(_03604_));
 sky130_fd_sc_hd__clkbuf_1 _17262_ (.A(_03604_),
    .X(_01566_));
 sky130_fd_sc_hd__buf_12 _17263_ (.A(_08958_),
    .X(_03605_));
 sky130_fd_sc_hd__nand2_8 _17264_ (.A(_06020_),
    .B(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__mux2_1 _17265_ (.A0(_03334_),
    .A1(net1775),
    .S(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__clkbuf_1 _17266_ (.A(_03607_),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _17267_ (.A0(_03337_),
    .A1(net906),
    .S(_03606_),
    .X(_03608_));
 sky130_fd_sc_hd__clkbuf_1 _17268_ (.A(_03608_),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _17269_ (.A0(_03339_),
    .A1(net1585),
    .S(_03606_),
    .X(_03609_));
 sky130_fd_sc_hd__clkbuf_1 _17270_ (.A(_03609_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _17271_ (.A0(_03341_),
    .A1(net1861),
    .S(_03606_),
    .X(_03610_));
 sky130_fd_sc_hd__clkbuf_1 _17272_ (.A(_03610_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _17273_ (.A0(_03343_),
    .A1(net984),
    .S(_03606_),
    .X(_03611_));
 sky130_fd_sc_hd__clkbuf_1 _17274_ (.A(_03611_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _17275_ (.A0(_03345_),
    .A1(net749),
    .S(_03606_),
    .X(_03612_));
 sky130_fd_sc_hd__clkbuf_1 _17276_ (.A(_03612_),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _17277_ (.A0(_03347_),
    .A1(net1556),
    .S(_03606_),
    .X(_03613_));
 sky130_fd_sc_hd__clkbuf_1 _17278_ (.A(_03613_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _17279_ (.A0(_03349_),
    .A1(net1649),
    .S(_03606_),
    .X(_03614_));
 sky130_fd_sc_hd__clkbuf_1 _17280_ (.A(_03614_),
    .X(_01574_));
 sky130_fd_sc_hd__nand2_8 _17281_ (.A(_06386_),
    .B(_03605_),
    .Y(_03615_));
 sky130_fd_sc_hd__mux2_1 _17282_ (.A0(_03334_),
    .A1(net857),
    .S(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__clkbuf_1 _17283_ (.A(_03616_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _17284_ (.A0(_03337_),
    .A1(net1063),
    .S(_03615_),
    .X(_03617_));
 sky130_fd_sc_hd__clkbuf_1 _17285_ (.A(_03617_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _17286_ (.A0(_03339_),
    .A1(net1469),
    .S(_03615_),
    .X(_03618_));
 sky130_fd_sc_hd__clkbuf_1 _17287_ (.A(_03618_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _17288_ (.A0(_03341_),
    .A1(net768),
    .S(_03615_),
    .X(_03619_));
 sky130_fd_sc_hd__clkbuf_1 _17289_ (.A(_03619_),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _17290_ (.A0(_03343_),
    .A1(net1264),
    .S(_03615_),
    .X(_03620_));
 sky130_fd_sc_hd__clkbuf_1 _17291_ (.A(_03620_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _17292_ (.A0(_03345_),
    .A1(net1042),
    .S(_03615_),
    .X(_03621_));
 sky130_fd_sc_hd__clkbuf_1 _17293_ (.A(_03621_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _17294_ (.A0(_03347_),
    .A1(net1252),
    .S(_03615_),
    .X(_03622_));
 sky130_fd_sc_hd__clkbuf_1 _17295_ (.A(_03622_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _17296_ (.A0(_03349_),
    .A1(net1389),
    .S(_03615_),
    .X(_03623_));
 sky130_fd_sc_hd__clkbuf_1 _17297_ (.A(_03623_),
    .X(_01582_));
 sky130_fd_sc_hd__and3_1 _17298_ (.A(_02266_),
    .B(_03595_),
    .C(_03516_),
    .X(_03624_));
 sky130_fd_sc_hd__buf_6 _17299_ (.A(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__mux2_1 _17300_ (.A0(net395),
    .A1(_03567_),
    .S(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__clkbuf_1 _17301_ (.A(_03626_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _17302_ (.A0(net1015),
    .A1(_03571_),
    .S(_03625_),
    .X(_03627_));
 sky130_fd_sc_hd__clkbuf_1 _17303_ (.A(_03627_),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _17304_ (.A0(net481),
    .A1(_03573_),
    .S(_03625_),
    .X(_03628_));
 sky130_fd_sc_hd__clkbuf_1 _17305_ (.A(_03628_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _17306_ (.A0(net340),
    .A1(_03575_),
    .S(_03625_),
    .X(_03629_));
 sky130_fd_sc_hd__clkbuf_1 _17307_ (.A(_03629_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _17308_ (.A0(net375),
    .A1(_03577_),
    .S(_03625_),
    .X(_03630_));
 sky130_fd_sc_hd__clkbuf_1 _17309_ (.A(_03630_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _17310_ (.A0(net540),
    .A1(_03579_),
    .S(_03625_),
    .X(_03631_));
 sky130_fd_sc_hd__clkbuf_1 _17311_ (.A(_03631_),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _17312_ (.A0(net1076),
    .A1(_03581_),
    .S(_03625_),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_1 _17313_ (.A(_03632_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _17314_ (.A0(net1292),
    .A1(_03583_),
    .S(_03625_),
    .X(_03633_));
 sky130_fd_sc_hd__clkbuf_1 _17315_ (.A(_03633_),
    .X(_01590_));
 sky130_fd_sc_hd__nand2_8 _17316_ (.A(_06217_),
    .B(_03605_),
    .Y(_03634_));
 sky130_fd_sc_hd__mux2_1 _17317_ (.A0(_03334_),
    .A1(net1479),
    .S(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__clkbuf_1 _17318_ (.A(_03635_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _17319_ (.A0(_03337_),
    .A1(net1052),
    .S(_03634_),
    .X(_03636_));
 sky130_fd_sc_hd__clkbuf_1 _17320_ (.A(_03636_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _17321_ (.A0(_03339_),
    .A1(net1484),
    .S(_03634_),
    .X(_03637_));
 sky130_fd_sc_hd__clkbuf_1 _17322_ (.A(_03637_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _17323_ (.A0(_03341_),
    .A1(net1366),
    .S(_03634_),
    .X(_03638_));
 sky130_fd_sc_hd__clkbuf_1 _17324_ (.A(_03638_),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _17325_ (.A0(_03343_),
    .A1(net1024),
    .S(_03634_),
    .X(_03639_));
 sky130_fd_sc_hd__clkbuf_1 _17326_ (.A(_03639_),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _17327_ (.A0(_03345_),
    .A1(net890),
    .S(_03634_),
    .X(_03640_));
 sky130_fd_sc_hd__clkbuf_1 _17328_ (.A(_03640_),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _17329_ (.A0(_03347_),
    .A1(net1273),
    .S(_03634_),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_1 _17330_ (.A(_03641_),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _17331_ (.A0(_03349_),
    .A1(net1784),
    .S(_03634_),
    .X(_03642_));
 sky130_fd_sc_hd__clkbuf_1 _17332_ (.A(_03642_),
    .X(_01598_));
 sky130_fd_sc_hd__and3_1 _17333_ (.A(_03595_),
    .B(_02286_),
    .C(_03516_),
    .X(_03643_));
 sky130_fd_sc_hd__buf_6 _17334_ (.A(_03643_),
    .X(_03644_));
 sky130_fd_sc_hd__mux2_1 _17335_ (.A0(net519),
    .A1(_03567_),
    .S(_03644_),
    .X(_03645_));
 sky130_fd_sc_hd__clkbuf_1 _17336_ (.A(_03645_),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _17337_ (.A0(net345),
    .A1(_03571_),
    .S(_03644_),
    .X(_03646_));
 sky130_fd_sc_hd__clkbuf_1 _17338_ (.A(_03646_),
    .X(_01600_));
 sky130_fd_sc_hd__mux2_1 _17339_ (.A0(net629),
    .A1(_03573_),
    .S(_03644_),
    .X(_03647_));
 sky130_fd_sc_hd__clkbuf_1 _17340_ (.A(_03647_),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _17341_ (.A0(net534),
    .A1(_03575_),
    .S(_03644_),
    .X(_03648_));
 sky130_fd_sc_hd__clkbuf_1 _17342_ (.A(_03648_),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_1 _17343_ (.A0(net523),
    .A1(_03577_),
    .S(_03644_),
    .X(_03649_));
 sky130_fd_sc_hd__clkbuf_1 _17344_ (.A(_03649_),
    .X(_01603_));
 sky130_fd_sc_hd__mux2_1 _17345_ (.A0(net661),
    .A1(_03579_),
    .S(_03644_),
    .X(_03650_));
 sky130_fd_sc_hd__clkbuf_1 _17346_ (.A(_03650_),
    .X(_01604_));
 sky130_fd_sc_hd__mux2_1 _17347_ (.A0(net855),
    .A1(_03581_),
    .S(_03644_),
    .X(_03651_));
 sky130_fd_sc_hd__clkbuf_1 _17348_ (.A(_03651_),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _17349_ (.A0(net1626),
    .A1(_03583_),
    .S(_03644_),
    .X(_03652_));
 sky130_fd_sc_hd__clkbuf_1 _17350_ (.A(_03652_),
    .X(_01606_));
 sky130_fd_sc_hd__and3_1 _17351_ (.A(_02297_),
    .B(_03595_),
    .C(_03516_),
    .X(_03653_));
 sky130_fd_sc_hd__clkbuf_8 _17352_ (.A(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__mux2_1 _17353_ (.A0(net875),
    .A1(_03567_),
    .S(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__clkbuf_1 _17354_ (.A(_03655_),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_1 _17355_ (.A0(net1651),
    .A1(_03571_),
    .S(_03654_),
    .X(_03656_));
 sky130_fd_sc_hd__clkbuf_1 _17356_ (.A(_03656_),
    .X(_01608_));
 sky130_fd_sc_hd__mux2_1 _17357_ (.A0(net851),
    .A1(_03573_),
    .S(_03654_),
    .X(_03657_));
 sky130_fd_sc_hd__clkbuf_1 _17358_ (.A(_03657_),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _17359_ (.A0(net869),
    .A1(_03575_),
    .S(_03654_),
    .X(_03658_));
 sky130_fd_sc_hd__clkbuf_1 _17360_ (.A(_03658_),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _17361_ (.A0(net564),
    .A1(_03577_),
    .S(_03654_),
    .X(_03659_));
 sky130_fd_sc_hd__clkbuf_1 _17362_ (.A(_03659_),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _17363_ (.A0(net431),
    .A1(_03579_),
    .S(_03654_),
    .X(_03660_));
 sky130_fd_sc_hd__clkbuf_1 _17364_ (.A(_03660_),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _17365_ (.A0(net1096),
    .A1(_03581_),
    .S(_03654_),
    .X(_03661_));
 sky130_fd_sc_hd__clkbuf_1 _17366_ (.A(_03661_),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _17367_ (.A0(net1073),
    .A1(_03583_),
    .S(_03654_),
    .X(_03662_));
 sky130_fd_sc_hd__clkbuf_1 _17368_ (.A(_03662_),
    .X(_01614_));
 sky130_fd_sc_hd__buf_2 _17369_ (.A(_08880_),
    .X(_03663_));
 sky130_fd_sc_hd__and3_1 _17370_ (.A(_03595_),
    .B(_06103_),
    .C(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__clkbuf_8 _17371_ (.A(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__mux2_1 _17372_ (.A0(net418),
    .A1(_03567_),
    .S(_03665_),
    .X(_03666_));
 sky130_fd_sc_hd__clkbuf_1 _17373_ (.A(_03666_),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _17374_ (.A0(net533),
    .A1(_03571_),
    .S(_03665_),
    .X(_03667_));
 sky130_fd_sc_hd__clkbuf_1 _17375_ (.A(_03667_),
    .X(_01616_));
 sky130_fd_sc_hd__mux2_1 _17376_ (.A0(net496),
    .A1(_03573_),
    .S(_03665_),
    .X(_03668_));
 sky130_fd_sc_hd__clkbuf_1 _17377_ (.A(_03668_),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _17378_ (.A0(net413),
    .A1(_03575_),
    .S(_03665_),
    .X(_03669_));
 sky130_fd_sc_hd__clkbuf_1 _17379_ (.A(_03669_),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_1 _17380_ (.A0(net651),
    .A1(_03577_),
    .S(_03665_),
    .X(_03670_));
 sky130_fd_sc_hd__clkbuf_1 _17381_ (.A(_03670_),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _17382_ (.A0(net326),
    .A1(_03579_),
    .S(_03665_),
    .X(_03671_));
 sky130_fd_sc_hd__clkbuf_1 _17383_ (.A(_03671_),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _17384_ (.A0(net467),
    .A1(_03581_),
    .S(_03665_),
    .X(_03672_));
 sky130_fd_sc_hd__clkbuf_1 _17385_ (.A(_03672_),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _17386_ (.A0(net944),
    .A1(_03583_),
    .S(_03665_),
    .X(_03673_));
 sky130_fd_sc_hd__clkbuf_1 _17387_ (.A(_03673_),
    .X(_01622_));
 sky130_fd_sc_hd__buf_6 _17388_ (.A(_09132_),
    .X(_03674_));
 sky130_fd_sc_hd__nand2_8 _17389_ (.A(_06479_),
    .B(_03605_),
    .Y(_03675_));
 sky130_fd_sc_hd__mux2_1 _17390_ (.A0(_03674_),
    .A1(\cur_mb_mem[184][0] ),
    .S(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__clkbuf_1 _17391_ (.A(_03676_),
    .X(_01623_));
 sky130_fd_sc_hd__buf_8 _17392_ (.A(_09136_),
    .X(_03677_));
 sky130_fd_sc_hd__mux2_1 _17393_ (.A0(_03677_),
    .A1(net1517),
    .S(_03675_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_1 _17394_ (.A(_03678_),
    .X(_01624_));
 sky130_fd_sc_hd__clkbuf_8 _17395_ (.A(_09139_),
    .X(_03679_));
 sky130_fd_sc_hd__mux2_1 _17396_ (.A0(_03679_),
    .A1(\cur_mb_mem[184][2] ),
    .S(_03675_),
    .X(_03680_));
 sky130_fd_sc_hd__clkbuf_1 _17397_ (.A(_03680_),
    .X(_01625_));
 sky130_fd_sc_hd__clkbuf_8 _17398_ (.A(_09142_),
    .X(_03681_));
 sky130_fd_sc_hd__mux2_1 _17399_ (.A0(_03681_),
    .A1(net681),
    .S(_03675_),
    .X(_03682_));
 sky130_fd_sc_hd__clkbuf_1 _17400_ (.A(_03682_),
    .X(_01626_));
 sky130_fd_sc_hd__clkbuf_8 _17401_ (.A(_09145_),
    .X(_03683_));
 sky130_fd_sc_hd__mux2_1 _17402_ (.A0(_03683_),
    .A1(net916),
    .S(_03675_),
    .X(_03684_));
 sky130_fd_sc_hd__clkbuf_1 _17403_ (.A(_03684_),
    .X(_01627_));
 sky130_fd_sc_hd__clkbuf_8 _17404_ (.A(_09148_),
    .X(_03685_));
 sky130_fd_sc_hd__mux2_1 _17405_ (.A0(_03685_),
    .A1(net953),
    .S(_03675_),
    .X(_03686_));
 sky130_fd_sc_hd__clkbuf_1 _17406_ (.A(_03686_),
    .X(_01628_));
 sky130_fd_sc_hd__buf_6 _17407_ (.A(_09151_),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_1 _17408_ (.A0(_03687_),
    .A1(net1579),
    .S(_03675_),
    .X(_03688_));
 sky130_fd_sc_hd__clkbuf_1 _17409_ (.A(_03688_),
    .X(_01629_));
 sky130_fd_sc_hd__buf_6 _17410_ (.A(_09154_),
    .X(_03689_));
 sky130_fd_sc_hd__mux2_1 _17411_ (.A0(_03689_),
    .A1(net1195),
    .S(_03675_),
    .X(_03690_));
 sky130_fd_sc_hd__clkbuf_1 _17412_ (.A(_03690_),
    .X(_01630_));
 sky130_fd_sc_hd__and3_1 _17413_ (.A(_08978_),
    .B(_03595_),
    .C(_03663_),
    .X(_03691_));
 sky130_fd_sc_hd__buf_4 _17414_ (.A(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__mux2_1 _17415_ (.A0(net1650),
    .A1(_03567_),
    .S(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__clkbuf_1 _17416_ (.A(_03693_),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_1 _17417_ (.A0(net1473),
    .A1(_03571_),
    .S(_03692_),
    .X(_03694_));
 sky130_fd_sc_hd__clkbuf_1 _17418_ (.A(_03694_),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_1 _17419_ (.A0(net1725),
    .A1(_03573_),
    .S(_03692_),
    .X(_03695_));
 sky130_fd_sc_hd__clkbuf_1 _17420_ (.A(_03695_),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _17421_ (.A0(net1751),
    .A1(_03575_),
    .S(_03692_),
    .X(_03696_));
 sky130_fd_sc_hd__clkbuf_1 _17422_ (.A(_03696_),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _17423_ (.A0(net700),
    .A1(_03577_),
    .S(_03692_),
    .X(_03697_));
 sky130_fd_sc_hd__clkbuf_1 _17424_ (.A(_03697_),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _17425_ (.A0(net514),
    .A1(_03579_),
    .S(_03692_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_1 _17426_ (.A(_03698_),
    .X(_01636_));
 sky130_fd_sc_hd__mux2_1 _17427_ (.A0(net1080),
    .A1(_03581_),
    .S(_03692_),
    .X(_03699_));
 sky130_fd_sc_hd__clkbuf_1 _17428_ (.A(_03699_),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _17429_ (.A0(net950),
    .A1(_03583_),
    .S(_03692_),
    .X(_03700_));
 sky130_fd_sc_hd__clkbuf_1 _17430_ (.A(_03700_),
    .X(_01638_));
 sky130_fd_sc_hd__and3_1 _17431_ (.A(_02353_),
    .B(_03595_),
    .C(_03663_),
    .X(_03701_));
 sky130_fd_sc_hd__clkbuf_8 _17432_ (.A(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__mux2_1 _17433_ (.A0(net604),
    .A1(_03567_),
    .S(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__clkbuf_1 _17434_ (.A(_03703_),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _17435_ (.A0(net521),
    .A1(_03571_),
    .S(_03702_),
    .X(_03704_));
 sky130_fd_sc_hd__clkbuf_1 _17436_ (.A(_03704_),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_1 _17437_ (.A0(net784),
    .A1(_03573_),
    .S(_03702_),
    .X(_03705_));
 sky130_fd_sc_hd__clkbuf_1 _17438_ (.A(_03705_),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _17439_ (.A0(net1630),
    .A1(_03575_),
    .S(_03702_),
    .X(_03706_));
 sky130_fd_sc_hd__clkbuf_1 _17440_ (.A(_03706_),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _17441_ (.A0(net492),
    .A1(_03577_),
    .S(_03702_),
    .X(_03707_));
 sky130_fd_sc_hd__clkbuf_1 _17442_ (.A(_03707_),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _17443_ (.A0(net430),
    .A1(_03579_),
    .S(_03702_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_1 _17444_ (.A(_03708_),
    .X(_01644_));
 sky130_fd_sc_hd__mux2_1 _17445_ (.A0(net1114),
    .A1(_03581_),
    .S(_03702_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_1 _17446_ (.A(_03709_),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _17447_ (.A0(net903),
    .A1(_03583_),
    .S(_03702_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_1 _17448_ (.A(_03710_),
    .X(_01646_));
 sky130_fd_sc_hd__and3_1 _17449_ (.A(_02526_),
    .B(_03595_),
    .C(_03663_),
    .X(_03711_));
 sky130_fd_sc_hd__buf_4 _17450_ (.A(_03711_),
    .X(_03712_));
 sky130_fd_sc_hd__mux2_1 _17451_ (.A0(net1231),
    .A1(_03567_),
    .S(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_1 _17452_ (.A(_03713_),
    .X(_01647_));
 sky130_fd_sc_hd__mux2_1 _17453_ (.A0(net929),
    .A1(_03571_),
    .S(_03712_),
    .X(_03714_));
 sky130_fd_sc_hd__clkbuf_1 _17454_ (.A(_03714_),
    .X(_01648_));
 sky130_fd_sc_hd__mux2_1 _17455_ (.A0(net753),
    .A1(_03573_),
    .S(_03712_),
    .X(_03715_));
 sky130_fd_sc_hd__clkbuf_1 _17456_ (.A(_03715_),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _17457_ (.A0(net412),
    .A1(_03575_),
    .S(_03712_),
    .X(_03716_));
 sky130_fd_sc_hd__clkbuf_1 _17458_ (.A(_03716_),
    .X(_01650_));
 sky130_fd_sc_hd__mux2_1 _17459_ (.A0(net370),
    .A1(_03577_),
    .S(_03712_),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_1 _17460_ (.A(_03717_),
    .X(_01651_));
 sky130_fd_sc_hd__mux2_1 _17461_ (.A0(net474),
    .A1(_03579_),
    .S(_03712_),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_1 _17462_ (.A(_03718_),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _17463_ (.A0(net476),
    .A1(_03581_),
    .S(_03712_),
    .X(_03719_));
 sky130_fd_sc_hd__clkbuf_1 _17464_ (.A(_03719_),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _17465_ (.A0(net878),
    .A1(_03583_),
    .S(_03712_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_1 _17466_ (.A(_03720_),
    .X(_01654_));
 sky130_fd_sc_hd__and3_1 _17467_ (.A(_02374_),
    .B(_03595_),
    .C(_03663_),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_8 _17468_ (.A(_03721_),
    .X(_03722_));
 sky130_fd_sc_hd__mux2_1 _17469_ (.A0(net312),
    .A1(_03567_),
    .S(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__clkbuf_1 _17470_ (.A(_03723_),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _17471_ (.A0(net516),
    .A1(_03571_),
    .S(_03722_),
    .X(_03724_));
 sky130_fd_sc_hd__clkbuf_1 _17472_ (.A(_03724_),
    .X(_01656_));
 sky130_fd_sc_hd__mux2_1 _17473_ (.A0(net1646),
    .A1(_03573_),
    .S(_03722_),
    .X(_03725_));
 sky130_fd_sc_hd__clkbuf_1 _17474_ (.A(_03725_),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _17475_ (.A0(net769),
    .A1(_03575_),
    .S(_03722_),
    .X(_03726_));
 sky130_fd_sc_hd__clkbuf_1 _17476_ (.A(_03726_),
    .X(_01658_));
 sky130_fd_sc_hd__mux2_1 _17477_ (.A0(net400),
    .A1(_03577_),
    .S(_03722_),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_1 _17478_ (.A(_03727_),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _17479_ (.A0(net319),
    .A1(_03579_),
    .S(_03722_),
    .X(_03728_));
 sky130_fd_sc_hd__clkbuf_1 _17480_ (.A(_03728_),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _17481_ (.A0(net323),
    .A1(_03581_),
    .S(_03722_),
    .X(_03729_));
 sky130_fd_sc_hd__clkbuf_1 _17482_ (.A(_03729_),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _17483_ (.A0(net353),
    .A1(_03583_),
    .S(_03722_),
    .X(_03730_));
 sky130_fd_sc_hd__clkbuf_1 _17484_ (.A(_03730_),
    .X(_01662_));
 sky130_fd_sc_hd__buf_4 _17485_ (.A(_08530_),
    .X(_03731_));
 sky130_fd_sc_hd__and3_1 _17486_ (.A(_09025_),
    .B(_06037_),
    .C(_03663_),
    .X(_03732_));
 sky130_fd_sc_hd__clkbuf_4 _17487_ (.A(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__mux2_1 _17488_ (.A0(\cur_mb_mem[189][0] ),
    .A1(_03731_),
    .S(_03733_),
    .X(_03734_));
 sky130_fd_sc_hd__clkbuf_1 _17489_ (.A(_03734_),
    .X(_01663_));
 sky130_fd_sc_hd__buf_4 _17490_ (.A(_08535_),
    .X(_03735_));
 sky130_fd_sc_hd__mux2_1 _17491_ (.A0(\cur_mb_mem[189][1] ),
    .A1(_03735_),
    .S(_03733_),
    .X(_03736_));
 sky130_fd_sc_hd__clkbuf_1 _17492_ (.A(_03736_),
    .X(_01664_));
 sky130_fd_sc_hd__buf_4 _17493_ (.A(_08538_),
    .X(_03737_));
 sky130_fd_sc_hd__mux2_1 _17494_ (.A0(\cur_mb_mem[189][2] ),
    .A1(_03737_),
    .S(_03733_),
    .X(_03738_));
 sky130_fd_sc_hd__clkbuf_1 _17495_ (.A(_03738_),
    .X(_01665_));
 sky130_fd_sc_hd__clkbuf_8 _17496_ (.A(_08541_),
    .X(_03739_));
 sky130_fd_sc_hd__mux2_1 _17497_ (.A0(\cur_mb_mem[189][3] ),
    .A1(_03739_),
    .S(_03733_),
    .X(_03740_));
 sky130_fd_sc_hd__clkbuf_1 _17498_ (.A(_03740_),
    .X(_01666_));
 sky130_fd_sc_hd__buf_4 _17499_ (.A(_08544_),
    .X(_03741_));
 sky130_fd_sc_hd__mux2_1 _17500_ (.A0(\cur_mb_mem[189][4] ),
    .A1(_03741_),
    .S(_03733_),
    .X(_03742_));
 sky130_fd_sc_hd__clkbuf_1 _17501_ (.A(_03742_),
    .X(_01667_));
 sky130_fd_sc_hd__buf_4 _17502_ (.A(_08547_),
    .X(_03743_));
 sky130_fd_sc_hd__mux2_1 _17503_ (.A0(\cur_mb_mem[189][5] ),
    .A1(_03743_),
    .S(_03733_),
    .X(_03744_));
 sky130_fd_sc_hd__clkbuf_1 _17504_ (.A(_03744_),
    .X(_01668_));
 sky130_fd_sc_hd__clkbuf_4 _17505_ (.A(_08550_),
    .X(_03745_));
 sky130_fd_sc_hd__mux2_1 _17506_ (.A0(\cur_mb_mem[189][6] ),
    .A1(_03745_),
    .S(_03733_),
    .X(_03746_));
 sky130_fd_sc_hd__clkbuf_1 _17507_ (.A(_03746_),
    .X(_01669_));
 sky130_fd_sc_hd__clkbuf_4 _17508_ (.A(_08553_),
    .X(_03747_));
 sky130_fd_sc_hd__mux2_1 _17509_ (.A0(\cur_mb_mem[189][7] ),
    .A1(_03747_),
    .S(_03733_),
    .X(_03748_));
 sky130_fd_sc_hd__clkbuf_1 _17510_ (.A(_03748_),
    .X(_01670_));
 sky130_fd_sc_hd__and3_1 _17511_ (.A(_03595_),
    .B(_06025_),
    .C(_03663_),
    .X(_03749_));
 sky130_fd_sc_hd__buf_4 _17512_ (.A(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__mux2_1 _17513_ (.A0(\cur_mb_mem[190][0] ),
    .A1(_03731_),
    .S(_03750_),
    .X(_03751_));
 sky130_fd_sc_hd__clkbuf_1 _17514_ (.A(_03751_),
    .X(_01671_));
 sky130_fd_sc_hd__mux2_1 _17515_ (.A0(\cur_mb_mem[190][1] ),
    .A1(_03735_),
    .S(_03750_),
    .X(_03752_));
 sky130_fd_sc_hd__clkbuf_1 _17516_ (.A(_03752_),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_1 _17517_ (.A0(\cur_mb_mem[190][2] ),
    .A1(_03737_),
    .S(_03750_),
    .X(_03753_));
 sky130_fd_sc_hd__clkbuf_1 _17518_ (.A(_03753_),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _17519_ (.A0(\cur_mb_mem[190][3] ),
    .A1(_03739_),
    .S(_03750_),
    .X(_03754_));
 sky130_fd_sc_hd__clkbuf_1 _17520_ (.A(_03754_),
    .X(_01674_));
 sky130_fd_sc_hd__mux2_1 _17521_ (.A0(\cur_mb_mem[190][4] ),
    .A1(_03741_),
    .S(_03750_),
    .X(_03755_));
 sky130_fd_sc_hd__clkbuf_1 _17522_ (.A(_03755_),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_1 _17523_ (.A0(\cur_mb_mem[190][5] ),
    .A1(_03743_),
    .S(_03750_),
    .X(_03756_));
 sky130_fd_sc_hd__clkbuf_1 _17524_ (.A(_03756_),
    .X(_01676_));
 sky130_fd_sc_hd__mux2_1 _17525_ (.A0(\cur_mb_mem[190][6] ),
    .A1(_03745_),
    .S(_03750_),
    .X(_03757_));
 sky130_fd_sc_hd__clkbuf_1 _17526_ (.A(_03757_),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _17527_ (.A0(\cur_mb_mem[190][7] ),
    .A1(_03747_),
    .S(_03750_),
    .X(_03758_));
 sky130_fd_sc_hd__clkbuf_1 _17528_ (.A(_03758_),
    .X(_01678_));
 sky130_fd_sc_hd__and3_1 _17529_ (.A(_02406_),
    .B(_06037_),
    .C(_03663_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_4 _17530_ (.A(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__mux2_1 _17531_ (.A0(\cur_mb_mem[191][0] ),
    .A1(_03731_),
    .S(_03760_),
    .X(_03761_));
 sky130_fd_sc_hd__clkbuf_1 _17532_ (.A(_03761_),
    .X(_01679_));
 sky130_fd_sc_hd__mux2_1 _17533_ (.A0(\cur_mb_mem[191][1] ),
    .A1(_03735_),
    .S(_03760_),
    .X(_03762_));
 sky130_fd_sc_hd__clkbuf_1 _17534_ (.A(_03762_),
    .X(_01680_));
 sky130_fd_sc_hd__mux2_1 _17535_ (.A0(\cur_mb_mem[191][2] ),
    .A1(_03737_),
    .S(_03760_),
    .X(_03763_));
 sky130_fd_sc_hd__clkbuf_1 _17536_ (.A(_03763_),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _17537_ (.A0(\cur_mb_mem[191][3] ),
    .A1(_03739_),
    .S(_03760_),
    .X(_03764_));
 sky130_fd_sc_hd__clkbuf_1 _17538_ (.A(_03764_),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _17539_ (.A0(\cur_mb_mem[191][4] ),
    .A1(_03741_),
    .S(_03760_),
    .X(_03765_));
 sky130_fd_sc_hd__clkbuf_1 _17540_ (.A(_03765_),
    .X(_01683_));
 sky130_fd_sc_hd__mux2_1 _17541_ (.A0(\cur_mb_mem[191][5] ),
    .A1(_03743_),
    .S(_03760_),
    .X(_03766_));
 sky130_fd_sc_hd__clkbuf_1 _17542_ (.A(_03766_),
    .X(_01684_));
 sky130_fd_sc_hd__mux2_1 _17543_ (.A0(\cur_mb_mem[191][6] ),
    .A1(_03745_),
    .S(_03760_),
    .X(_03767_));
 sky130_fd_sc_hd__clkbuf_1 _17544_ (.A(_03767_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _17545_ (.A0(\cur_mb_mem[191][7] ),
    .A1(_03747_),
    .S(_03760_),
    .X(_03768_));
 sky130_fd_sc_hd__clkbuf_1 _17546_ (.A(_03768_),
    .X(_01686_));
 sky130_fd_sc_hd__buf_4 _17547_ (.A(_06094_),
    .X(_03769_));
 sky130_fd_sc_hd__nand2_8 _17548_ (.A(_03769_),
    .B(_08882_),
    .Y(_03770_));
 sky130_fd_sc_hd__mux2_1 _17549_ (.A0(_03674_),
    .A1(net1443),
    .S(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__clkbuf_1 _17550_ (.A(_03771_),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _17551_ (.A0(_03677_),
    .A1(net808),
    .S(_03770_),
    .X(_03772_));
 sky130_fd_sc_hd__clkbuf_1 _17552_ (.A(_03772_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _17553_ (.A0(_03679_),
    .A1(net941),
    .S(_03770_),
    .X(_03773_));
 sky130_fd_sc_hd__clkbuf_1 _17554_ (.A(_03773_),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_1 _17555_ (.A0(_03681_),
    .A1(net1392),
    .S(_03770_),
    .X(_03774_));
 sky130_fd_sc_hd__clkbuf_1 _17556_ (.A(_03774_),
    .X(_01690_));
 sky130_fd_sc_hd__mux2_1 _17557_ (.A0(_03683_),
    .A1(net1606),
    .S(_03770_),
    .X(_03775_));
 sky130_fd_sc_hd__clkbuf_1 _17558_ (.A(_03775_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _17559_ (.A0(_03685_),
    .A1(net1048),
    .S(_03770_),
    .X(_03776_));
 sky130_fd_sc_hd__clkbuf_1 _17560_ (.A(_03776_),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_1 _17561_ (.A0(_03687_),
    .A1(net1045),
    .S(_03770_),
    .X(_03777_));
 sky130_fd_sc_hd__clkbuf_1 _17562_ (.A(_03777_),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _17563_ (.A0(_03689_),
    .A1(net636),
    .S(_03770_),
    .X(_03778_));
 sky130_fd_sc_hd__clkbuf_1 _17564_ (.A(_03778_),
    .X(_01694_));
 sky130_fd_sc_hd__nand2_8 _17565_ (.A(_06354_),
    .B(_03605_),
    .Y(_03779_));
 sky130_fd_sc_hd__mux2_1 _17566_ (.A0(_03674_),
    .A1(net794),
    .S(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__clkbuf_1 _17567_ (.A(_03780_),
    .X(_01695_));
 sky130_fd_sc_hd__mux2_1 _17568_ (.A0(_03677_),
    .A1(net1713),
    .S(_03779_),
    .X(_03781_));
 sky130_fd_sc_hd__clkbuf_1 _17569_ (.A(_03781_),
    .X(_01696_));
 sky130_fd_sc_hd__mux2_1 _17570_ (.A0(_03679_),
    .A1(net1279),
    .S(_03779_),
    .X(_03782_));
 sky130_fd_sc_hd__clkbuf_1 _17571_ (.A(_03782_),
    .X(_01697_));
 sky130_fd_sc_hd__mux2_1 _17572_ (.A0(_03681_),
    .A1(net396),
    .S(_03779_),
    .X(_03783_));
 sky130_fd_sc_hd__clkbuf_1 _17573_ (.A(_03783_),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _17574_ (.A0(_03683_),
    .A1(net1126),
    .S(_03779_),
    .X(_03784_));
 sky130_fd_sc_hd__clkbuf_1 _17575_ (.A(_03784_),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _17576_ (.A0(_03685_),
    .A1(net1553),
    .S(_03779_),
    .X(_03785_));
 sky130_fd_sc_hd__clkbuf_1 _17577_ (.A(_03785_),
    .X(_01700_));
 sky130_fd_sc_hd__mux2_1 _17578_ (.A0(_03687_),
    .A1(net1161),
    .S(_03779_),
    .X(_03786_));
 sky130_fd_sc_hd__clkbuf_1 _17579_ (.A(_03786_),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_1 _17580_ (.A0(_03689_),
    .A1(net1320),
    .S(_03779_),
    .X(_03787_));
 sky130_fd_sc_hd__clkbuf_1 _17581_ (.A(_03787_),
    .X(_01702_));
 sky130_fd_sc_hd__nand2_8 _17582_ (.A(_06083_),
    .B(_03605_),
    .Y(_03788_));
 sky130_fd_sc_hd__mux2_1 _17583_ (.A0(_03674_),
    .A1(net498),
    .S(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__clkbuf_1 _17584_ (.A(_03789_),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _17585_ (.A0(_03677_),
    .A1(net1265),
    .S(_03788_),
    .X(_03790_));
 sky130_fd_sc_hd__clkbuf_1 _17586_ (.A(_03790_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _17587_ (.A0(_03679_),
    .A1(net1170),
    .S(_03788_),
    .X(_03791_));
 sky130_fd_sc_hd__clkbuf_1 _17588_ (.A(_03791_),
    .X(_01705_));
 sky130_fd_sc_hd__mux2_1 _17589_ (.A0(_03681_),
    .A1(net719),
    .S(_03788_),
    .X(_03792_));
 sky130_fd_sc_hd__clkbuf_1 _17590_ (.A(_03792_),
    .X(_01706_));
 sky130_fd_sc_hd__mux2_1 _17591_ (.A0(_03683_),
    .A1(net977),
    .S(_03788_),
    .X(_03793_));
 sky130_fd_sc_hd__clkbuf_1 _17592_ (.A(_03793_),
    .X(_01707_));
 sky130_fd_sc_hd__mux2_1 _17593_ (.A0(_03685_),
    .A1(net1147),
    .S(_03788_),
    .X(_03794_));
 sky130_fd_sc_hd__clkbuf_1 _17594_ (.A(_03794_),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_1 _17595_ (.A0(_03687_),
    .A1(net1388),
    .S(_03788_),
    .X(_03795_));
 sky130_fd_sc_hd__clkbuf_1 _17596_ (.A(_03795_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _17597_ (.A0(_03689_),
    .A1(net1070),
    .S(_03788_),
    .X(_03796_));
 sky130_fd_sc_hd__clkbuf_1 _17598_ (.A(_03796_),
    .X(_01710_));
 sky130_fd_sc_hd__and3_1 _17599_ (.A(_02266_),
    .B(_03769_),
    .C(_03663_),
    .X(_03797_));
 sky130_fd_sc_hd__buf_4 _17600_ (.A(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__mux2_1 _17601_ (.A0(\cur_mb_mem[195][0] ),
    .A1(_03731_),
    .S(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__clkbuf_1 _17602_ (.A(_03799_),
    .X(_01711_));
 sky130_fd_sc_hd__mux2_1 _17603_ (.A0(\cur_mb_mem[195][1] ),
    .A1(_03735_),
    .S(_03798_),
    .X(_03800_));
 sky130_fd_sc_hd__clkbuf_1 _17604_ (.A(_03800_),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _17605_ (.A0(\cur_mb_mem[195][2] ),
    .A1(_03737_),
    .S(_03798_),
    .X(_03801_));
 sky130_fd_sc_hd__clkbuf_1 _17606_ (.A(_03801_),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _17607_ (.A0(\cur_mb_mem[195][3] ),
    .A1(_03739_),
    .S(_03798_),
    .X(_03802_));
 sky130_fd_sc_hd__clkbuf_1 _17608_ (.A(_03802_),
    .X(_01714_));
 sky130_fd_sc_hd__mux2_1 _17609_ (.A0(net1877),
    .A1(_03741_),
    .S(_03798_),
    .X(_03803_));
 sky130_fd_sc_hd__clkbuf_1 _17610_ (.A(_03803_),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_1 _17611_ (.A0(net1872),
    .A1(_03743_),
    .S(_03798_),
    .X(_03804_));
 sky130_fd_sc_hd__clkbuf_1 _17612_ (.A(_03804_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _17613_ (.A0(\cur_mb_mem[195][6] ),
    .A1(_03745_),
    .S(_03798_),
    .X(_03805_));
 sky130_fd_sc_hd__clkbuf_1 _17614_ (.A(_03805_),
    .X(_01717_));
 sky130_fd_sc_hd__mux2_1 _17615_ (.A0(\cur_mb_mem[195][7] ),
    .A1(_03747_),
    .S(_03798_),
    .X(_03806_));
 sky130_fd_sc_hd__clkbuf_1 _17616_ (.A(_03806_),
    .X(_01718_));
 sky130_fd_sc_hd__nand3_4 _17617_ (.A(_06223_),
    .B(_03769_),
    .C(_08901_),
    .Y(_03807_));
 sky130_fd_sc_hd__mux2_1 _17618_ (.A0(_03674_),
    .A1(net1182),
    .S(_03807_),
    .X(_03808_));
 sky130_fd_sc_hd__clkbuf_1 _17619_ (.A(_03808_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _17620_ (.A0(_03677_),
    .A1(net575),
    .S(net214),
    .X(_03809_));
 sky130_fd_sc_hd__clkbuf_1 _17621_ (.A(_03809_),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _17622_ (.A0(_03679_),
    .A1(net722),
    .S(net214),
    .X(_03810_));
 sky130_fd_sc_hd__clkbuf_1 _17623_ (.A(_03810_),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _17624_ (.A0(_03681_),
    .A1(net1300),
    .S(_03807_),
    .X(_03811_));
 sky130_fd_sc_hd__clkbuf_1 _17625_ (.A(_03811_),
    .X(_01722_));
 sky130_fd_sc_hd__mux2_1 _17626_ (.A0(_03683_),
    .A1(net536),
    .S(_03807_),
    .X(_03812_));
 sky130_fd_sc_hd__clkbuf_1 _17627_ (.A(_03812_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _17628_ (.A0(_03685_),
    .A1(net721),
    .S(_03807_),
    .X(_03813_));
 sky130_fd_sc_hd__clkbuf_1 _17629_ (.A(_03813_),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _17630_ (.A0(_03687_),
    .A1(net1548),
    .S(net214),
    .X(_03814_));
 sky130_fd_sc_hd__clkbuf_1 _17631_ (.A(_03814_),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_1 _17632_ (.A0(_03689_),
    .A1(net1741),
    .S(net214),
    .X(_03815_));
 sky130_fd_sc_hd__clkbuf_1 _17633_ (.A(_03815_),
    .X(_01726_));
 sky130_fd_sc_hd__and3_1 _17634_ (.A(_03769_),
    .B(_02286_),
    .C(_03663_),
    .X(_03816_));
 sky130_fd_sc_hd__buf_4 _17635_ (.A(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__mux2_1 _17636_ (.A0(\cur_mb_mem[197][0] ),
    .A1(_03731_),
    .S(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__clkbuf_1 _17637_ (.A(_03818_),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _17638_ (.A0(\cur_mb_mem[197][1] ),
    .A1(_03735_),
    .S(_03817_),
    .X(_03819_));
 sky130_fd_sc_hd__clkbuf_1 _17639_ (.A(_03819_),
    .X(_01728_));
 sky130_fd_sc_hd__mux2_1 _17640_ (.A0(\cur_mb_mem[197][2] ),
    .A1(_03737_),
    .S(_03817_),
    .X(_03820_));
 sky130_fd_sc_hd__clkbuf_1 _17641_ (.A(_03820_),
    .X(_01729_));
 sky130_fd_sc_hd__mux2_1 _17642_ (.A0(\cur_mb_mem[197][3] ),
    .A1(_03739_),
    .S(_03817_),
    .X(_03821_));
 sky130_fd_sc_hd__clkbuf_1 _17643_ (.A(_03821_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _17644_ (.A0(net1993),
    .A1(_03741_),
    .S(_03817_),
    .X(_03822_));
 sky130_fd_sc_hd__clkbuf_1 _17645_ (.A(_03822_),
    .X(_01731_));
 sky130_fd_sc_hd__mux2_1 _17646_ (.A0(net1985),
    .A1(_03743_),
    .S(_03817_),
    .X(_03823_));
 sky130_fd_sc_hd__clkbuf_1 _17647_ (.A(_03823_),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_1 _17648_ (.A0(\cur_mb_mem[197][6] ),
    .A1(_03745_),
    .S(_03817_),
    .X(_03824_));
 sky130_fd_sc_hd__clkbuf_1 _17649_ (.A(_03824_),
    .X(_01733_));
 sky130_fd_sc_hd__mux2_1 _17650_ (.A0(\cur_mb_mem[197][7] ),
    .A1(_03747_),
    .S(_03817_),
    .X(_03825_));
 sky130_fd_sc_hd__clkbuf_1 _17651_ (.A(_03825_),
    .X(_01734_));
 sky130_fd_sc_hd__clkbuf_2 _17652_ (.A(_08880_),
    .X(_03826_));
 sky130_fd_sc_hd__and3_1 _17653_ (.A(_02297_),
    .B(_03769_),
    .C(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__buf_4 _17654_ (.A(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__mux2_1 _17655_ (.A0(net1945),
    .A1(_03731_),
    .S(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__clkbuf_1 _17656_ (.A(_03829_),
    .X(_01735_));
 sky130_fd_sc_hd__mux2_1 _17657_ (.A0(\cur_mb_mem[198][1] ),
    .A1(_03735_),
    .S(_03828_),
    .X(_03830_));
 sky130_fd_sc_hd__clkbuf_1 _17658_ (.A(_03830_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _17659_ (.A0(\cur_mb_mem[198][2] ),
    .A1(_03737_),
    .S(_03828_),
    .X(_03831_));
 sky130_fd_sc_hd__clkbuf_1 _17660_ (.A(_03831_),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _17661_ (.A0(\cur_mb_mem[198][3] ),
    .A1(_03739_),
    .S(_03828_),
    .X(_03832_));
 sky130_fd_sc_hd__clkbuf_1 _17662_ (.A(_03832_),
    .X(_01738_));
 sky130_fd_sc_hd__mux2_1 _17663_ (.A0(\cur_mb_mem[198][4] ),
    .A1(_03741_),
    .S(_03828_),
    .X(_03833_));
 sky130_fd_sc_hd__clkbuf_1 _17664_ (.A(_03833_),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _17665_ (.A0(net1981),
    .A1(_03743_),
    .S(_03828_),
    .X(_03834_));
 sky130_fd_sc_hd__clkbuf_1 _17666_ (.A(_03834_),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _17667_ (.A0(\cur_mb_mem[198][6] ),
    .A1(_03745_),
    .S(_03828_),
    .X(_03835_));
 sky130_fd_sc_hd__clkbuf_1 _17668_ (.A(_03835_),
    .X(_01741_));
 sky130_fd_sc_hd__mux2_1 _17669_ (.A0(\cur_mb_mem[198][7] ),
    .A1(_03747_),
    .S(_03828_),
    .X(_03836_));
 sky130_fd_sc_hd__clkbuf_1 _17670_ (.A(_03836_),
    .X(_01742_));
 sky130_fd_sc_hd__and3_1 _17671_ (.A(_03769_),
    .B(_06103_),
    .C(_03826_),
    .X(_03837_));
 sky130_fd_sc_hd__buf_4 _17672_ (.A(_03837_),
    .X(_03838_));
 sky130_fd_sc_hd__mux2_1 _17673_ (.A0(\cur_mb_mem[199][0] ),
    .A1(_03731_),
    .S(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__clkbuf_1 _17674_ (.A(_03839_),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _17675_ (.A0(\cur_mb_mem[199][1] ),
    .A1(_03735_),
    .S(_03838_),
    .X(_03840_));
 sky130_fd_sc_hd__clkbuf_1 _17676_ (.A(_03840_),
    .X(_01744_));
 sky130_fd_sc_hd__mux2_1 _17677_ (.A0(\cur_mb_mem[199][2] ),
    .A1(_03737_),
    .S(_03838_),
    .X(_03841_));
 sky130_fd_sc_hd__clkbuf_1 _17678_ (.A(_03841_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_1 _17679_ (.A0(\cur_mb_mem[199][3] ),
    .A1(_03739_),
    .S(_03838_),
    .X(_03842_));
 sky130_fd_sc_hd__clkbuf_1 _17680_ (.A(_03842_),
    .X(_01746_));
 sky130_fd_sc_hd__mux2_1 _17681_ (.A0(\cur_mb_mem[199][4] ),
    .A1(_03741_),
    .S(_03838_),
    .X(_03843_));
 sky130_fd_sc_hd__clkbuf_1 _17682_ (.A(_03843_),
    .X(_01747_));
 sky130_fd_sc_hd__mux2_1 _17683_ (.A0(\cur_mb_mem[199][5] ),
    .A1(_03743_),
    .S(_03838_),
    .X(_03844_));
 sky130_fd_sc_hd__clkbuf_1 _17684_ (.A(_03844_),
    .X(_01748_));
 sky130_fd_sc_hd__mux2_1 _17685_ (.A0(\cur_mb_mem[199][6] ),
    .A1(_03745_),
    .S(_03838_),
    .X(_03845_));
 sky130_fd_sc_hd__clkbuf_1 _17686_ (.A(_03845_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _17687_ (.A0(\cur_mb_mem[199][7] ),
    .A1(_03747_),
    .S(_03838_),
    .X(_03846_));
 sky130_fd_sc_hd__clkbuf_1 _17688_ (.A(_03846_),
    .X(_01750_));
 sky130_fd_sc_hd__nand2_8 _17689_ (.A(_06457_),
    .B(_03605_),
    .Y(_03847_));
 sky130_fd_sc_hd__mux2_1 _17690_ (.A0(_03674_),
    .A1(net667),
    .S(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__clkbuf_1 _17691_ (.A(_03848_),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _17692_ (.A0(_03677_),
    .A1(net1435),
    .S(_03847_),
    .X(_03849_));
 sky130_fd_sc_hd__clkbuf_1 _17693_ (.A(_03849_),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _17694_ (.A0(_03679_),
    .A1(net730),
    .S(_03847_),
    .X(_03850_));
 sky130_fd_sc_hd__clkbuf_1 _17695_ (.A(_03850_),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _17696_ (.A0(_03681_),
    .A1(net1764),
    .S(_03847_),
    .X(_03851_));
 sky130_fd_sc_hd__clkbuf_1 _17697_ (.A(_03851_),
    .X(_01754_));
 sky130_fd_sc_hd__mux2_1 _17698_ (.A0(_03683_),
    .A1(net1284),
    .S(_03847_),
    .X(_03852_));
 sky130_fd_sc_hd__clkbuf_1 _17699_ (.A(_03852_),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_1 _17700_ (.A0(_03685_),
    .A1(net1797),
    .S(_03847_),
    .X(_03853_));
 sky130_fd_sc_hd__clkbuf_1 _17701_ (.A(_03853_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _17702_ (.A0(_03687_),
    .A1(net1427),
    .S(_03847_),
    .X(_03854_));
 sky130_fd_sc_hd__clkbuf_1 _17703_ (.A(_03854_),
    .X(_01757_));
 sky130_fd_sc_hd__mux2_1 _17704_ (.A0(_03689_),
    .A1(net1472),
    .S(_03847_),
    .X(_03855_));
 sky130_fd_sc_hd__clkbuf_1 _17705_ (.A(_03855_),
    .X(_01758_));
 sky130_fd_sc_hd__and3_1 _17706_ (.A(_08978_),
    .B(_03769_),
    .C(_03826_),
    .X(_03856_));
 sky130_fd_sc_hd__buf_4 _17707_ (.A(_03856_),
    .X(_03857_));
 sky130_fd_sc_hd__mux2_1 _17708_ (.A0(\cur_mb_mem[201][0] ),
    .A1(_03731_),
    .S(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__clkbuf_1 _17709_ (.A(_03858_),
    .X(_01759_));
 sky130_fd_sc_hd__mux2_1 _17710_ (.A0(\cur_mb_mem[201][1] ),
    .A1(_03735_),
    .S(_03857_),
    .X(_03859_));
 sky130_fd_sc_hd__clkbuf_1 _17711_ (.A(_03859_),
    .X(_01760_));
 sky130_fd_sc_hd__mux2_1 _17712_ (.A0(\cur_mb_mem[201][2] ),
    .A1(_03737_),
    .S(_03857_),
    .X(_03860_));
 sky130_fd_sc_hd__clkbuf_1 _17713_ (.A(_03860_),
    .X(_01761_));
 sky130_fd_sc_hd__mux2_1 _17714_ (.A0(\cur_mb_mem[201][3] ),
    .A1(_03739_),
    .S(_03857_),
    .X(_03861_));
 sky130_fd_sc_hd__clkbuf_1 _17715_ (.A(_03861_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _17716_ (.A0(net1883),
    .A1(_03741_),
    .S(_03857_),
    .X(_03862_));
 sky130_fd_sc_hd__clkbuf_1 _17717_ (.A(_03862_),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _17718_ (.A0(net1923),
    .A1(_03743_),
    .S(_03857_),
    .X(_03863_));
 sky130_fd_sc_hd__clkbuf_1 _17719_ (.A(_03863_),
    .X(_01764_));
 sky130_fd_sc_hd__mux2_1 _17720_ (.A0(\cur_mb_mem[201][6] ),
    .A1(_03745_),
    .S(_03857_),
    .X(_03864_));
 sky130_fd_sc_hd__clkbuf_1 _17721_ (.A(_03864_),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _17722_ (.A0(\cur_mb_mem[201][7] ),
    .A1(_03747_),
    .S(_03857_),
    .X(_03865_));
 sky130_fd_sc_hd__clkbuf_1 _17723_ (.A(_03865_),
    .X(_01766_));
 sky130_fd_sc_hd__and3_1 _17724_ (.A(_02353_),
    .B(_03769_),
    .C(_03826_),
    .X(_03866_));
 sky130_fd_sc_hd__clkbuf_4 _17725_ (.A(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__mux2_1 _17726_ (.A0(\cur_mb_mem[202][0] ),
    .A1(_03731_),
    .S(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__clkbuf_1 _17727_ (.A(_03868_),
    .X(_01767_));
 sky130_fd_sc_hd__mux2_1 _17728_ (.A0(\cur_mb_mem[202][1] ),
    .A1(_03735_),
    .S(_03867_),
    .X(_03869_));
 sky130_fd_sc_hd__clkbuf_1 _17729_ (.A(_03869_),
    .X(_01768_));
 sky130_fd_sc_hd__mux2_1 _17730_ (.A0(net1958),
    .A1(_03737_),
    .S(_03867_),
    .X(_03870_));
 sky130_fd_sc_hd__clkbuf_1 _17731_ (.A(_03870_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _17732_ (.A0(\cur_mb_mem[202][3] ),
    .A1(_03739_),
    .S(_03867_),
    .X(_03871_));
 sky130_fd_sc_hd__clkbuf_1 _17733_ (.A(_03871_),
    .X(_01770_));
 sky130_fd_sc_hd__mux2_1 _17734_ (.A0(net1966),
    .A1(_03741_),
    .S(_03867_),
    .X(_03872_));
 sky130_fd_sc_hd__clkbuf_1 _17735_ (.A(_03872_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _17736_ (.A0(\cur_mb_mem[202][5] ),
    .A1(_03743_),
    .S(_03867_),
    .X(_03873_));
 sky130_fd_sc_hd__clkbuf_1 _17737_ (.A(_03873_),
    .X(_01772_));
 sky130_fd_sc_hd__mux2_1 _17738_ (.A0(\cur_mb_mem[202][6] ),
    .A1(_03745_),
    .S(_03867_),
    .X(_03874_));
 sky130_fd_sc_hd__clkbuf_1 _17739_ (.A(_03874_),
    .X(_01773_));
 sky130_fd_sc_hd__mux2_1 _17740_ (.A0(\cur_mb_mem[202][7] ),
    .A1(_03747_),
    .S(_03867_),
    .X(_03875_));
 sky130_fd_sc_hd__clkbuf_1 _17741_ (.A(_03875_),
    .X(_01774_));
 sky130_fd_sc_hd__and3_1 _17742_ (.A(_02526_),
    .B(_03769_),
    .C(_03826_),
    .X(_03876_));
 sky130_fd_sc_hd__clkbuf_4 _17743_ (.A(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__mux2_1 _17744_ (.A0(\cur_mb_mem[203][0] ),
    .A1(_03731_),
    .S(_03877_),
    .X(_03878_));
 sky130_fd_sc_hd__clkbuf_1 _17745_ (.A(_03878_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _17746_ (.A0(\cur_mb_mem[203][1] ),
    .A1(_03735_),
    .S(_03877_),
    .X(_03879_));
 sky130_fd_sc_hd__clkbuf_1 _17747_ (.A(_03879_),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _17748_ (.A0(\cur_mb_mem[203][2] ),
    .A1(_03737_),
    .S(_03877_),
    .X(_03880_));
 sky130_fd_sc_hd__clkbuf_1 _17749_ (.A(_03880_),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_1 _17750_ (.A0(\cur_mb_mem[203][3] ),
    .A1(_03739_),
    .S(_03877_),
    .X(_03881_));
 sky130_fd_sc_hd__clkbuf_1 _17751_ (.A(_03881_),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _17752_ (.A0(net1977),
    .A1(_03741_),
    .S(_03877_),
    .X(_03882_));
 sky130_fd_sc_hd__clkbuf_1 _17753_ (.A(_03882_),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _17754_ (.A0(\cur_mb_mem[203][5] ),
    .A1(_03743_),
    .S(_03877_),
    .X(_03883_));
 sky130_fd_sc_hd__clkbuf_1 _17755_ (.A(_03883_),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _17756_ (.A0(\cur_mb_mem[203][6] ),
    .A1(_03745_),
    .S(_03877_),
    .X(_03884_));
 sky130_fd_sc_hd__clkbuf_1 _17757_ (.A(_03884_),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _17758_ (.A0(\cur_mb_mem[203][7] ),
    .A1(_03747_),
    .S(_03877_),
    .X(_03885_));
 sky130_fd_sc_hd__clkbuf_1 _17759_ (.A(_03885_),
    .X(_01782_));
 sky130_fd_sc_hd__buf_4 _17760_ (.A(_08530_),
    .X(_03886_));
 sky130_fd_sc_hd__and3_1 _17761_ (.A(_02374_),
    .B(_03769_),
    .C(_03826_),
    .X(_03887_));
 sky130_fd_sc_hd__buf_4 _17762_ (.A(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__mux2_1 _17763_ (.A0(net1991),
    .A1(_03886_),
    .S(_03888_),
    .X(_03889_));
 sky130_fd_sc_hd__clkbuf_1 _17764_ (.A(_03889_),
    .X(_01783_));
 sky130_fd_sc_hd__clkbuf_4 _17765_ (.A(_08535_),
    .X(_03890_));
 sky130_fd_sc_hd__mux2_1 _17766_ (.A0(\cur_mb_mem[204][1] ),
    .A1(_03890_),
    .S(_03888_),
    .X(_03891_));
 sky130_fd_sc_hd__clkbuf_1 _17767_ (.A(_03891_),
    .X(_01784_));
 sky130_fd_sc_hd__buf_4 _17768_ (.A(_08538_),
    .X(_03892_));
 sky130_fd_sc_hd__mux2_1 _17769_ (.A0(\cur_mb_mem[204][2] ),
    .A1(_03892_),
    .S(_03888_),
    .X(_03893_));
 sky130_fd_sc_hd__clkbuf_1 _17770_ (.A(_03893_),
    .X(_01785_));
 sky130_fd_sc_hd__buf_4 _17771_ (.A(_08541_),
    .X(_03894_));
 sky130_fd_sc_hd__mux2_1 _17772_ (.A0(\cur_mb_mem[204][3] ),
    .A1(_03894_),
    .S(_03888_),
    .X(_03895_));
 sky130_fd_sc_hd__clkbuf_1 _17773_ (.A(_03895_),
    .X(_01786_));
 sky130_fd_sc_hd__clkbuf_4 _17774_ (.A(_08544_),
    .X(_03896_));
 sky130_fd_sc_hd__mux2_1 _17775_ (.A0(net1740),
    .A1(_03896_),
    .S(_03888_),
    .X(_03897_));
 sky130_fd_sc_hd__clkbuf_1 _17776_ (.A(_03897_),
    .X(_01787_));
 sky130_fd_sc_hd__buf_4 _17777_ (.A(_08547_),
    .X(_03898_));
 sky130_fd_sc_hd__mux2_1 _17778_ (.A0(net1804),
    .A1(_03898_),
    .S(_03888_),
    .X(_03899_));
 sky130_fd_sc_hd__clkbuf_1 _17779_ (.A(_03899_),
    .X(_01788_));
 sky130_fd_sc_hd__clkbuf_4 _17780_ (.A(_08550_),
    .X(_03900_));
 sky130_fd_sc_hd__mux2_1 _17781_ (.A0(net1964),
    .A1(_03900_),
    .S(_03888_),
    .X(_03901_));
 sky130_fd_sc_hd__clkbuf_1 _17782_ (.A(_03901_),
    .X(_01789_));
 sky130_fd_sc_hd__clkbuf_4 _17783_ (.A(_08553_),
    .X(_03902_));
 sky130_fd_sc_hd__mux2_1 _17784_ (.A0(\cur_mb_mem[204][7] ),
    .A1(_03902_),
    .S(_03888_),
    .X(_03903_));
 sky130_fd_sc_hd__clkbuf_1 _17785_ (.A(_03903_),
    .X(_01790_));
 sky130_fd_sc_hd__and3_1 _17786_ (.A(_09025_),
    .B(_06094_),
    .C(_03826_),
    .X(_03904_));
 sky130_fd_sc_hd__clkbuf_4 _17787_ (.A(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__mux2_1 _17788_ (.A0(\cur_mb_mem[205][0] ),
    .A1(_03886_),
    .S(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__clkbuf_1 _17789_ (.A(_03906_),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _17790_ (.A0(net1769),
    .A1(_03890_),
    .S(_03905_),
    .X(_03907_));
 sky130_fd_sc_hd__clkbuf_1 _17791_ (.A(_03907_),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _17792_ (.A0(net1634),
    .A1(_03892_),
    .S(_03905_),
    .X(_03908_));
 sky130_fd_sc_hd__clkbuf_1 _17793_ (.A(_03908_),
    .X(_01793_));
 sky130_fd_sc_hd__mux2_1 _17794_ (.A0(\cur_mb_mem[205][3] ),
    .A1(_03894_),
    .S(_03905_),
    .X(_03909_));
 sky130_fd_sc_hd__clkbuf_1 _17795_ (.A(_03909_),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_1 _17796_ (.A0(net1628),
    .A1(_03896_),
    .S(_03905_),
    .X(_03910_));
 sky130_fd_sc_hd__clkbuf_1 _17797_ (.A(_03910_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _17798_ (.A0(net1676),
    .A1(_03898_),
    .S(_03905_),
    .X(_03911_));
 sky130_fd_sc_hd__clkbuf_1 _17799_ (.A(_03911_),
    .X(_01796_));
 sky130_fd_sc_hd__mux2_1 _17800_ (.A0(\cur_mb_mem[205][6] ),
    .A1(_03900_),
    .S(_03905_),
    .X(_03912_));
 sky130_fd_sc_hd__clkbuf_1 _17801_ (.A(_03912_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _17802_ (.A0(\cur_mb_mem[205][7] ),
    .A1(_03902_),
    .S(_03905_),
    .X(_03913_));
 sky130_fd_sc_hd__clkbuf_1 _17803_ (.A(_03913_),
    .X(_01798_));
 sky130_fd_sc_hd__and3_1 _17804_ (.A(_09036_),
    .B(_06094_),
    .C(_03826_),
    .X(_03914_));
 sky130_fd_sc_hd__buf_4 _17805_ (.A(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__mux2_1 _17806_ (.A0(\cur_mb_mem[206][0] ),
    .A1(_03886_),
    .S(_03915_),
    .X(_03916_));
 sky130_fd_sc_hd__clkbuf_1 _17807_ (.A(_03916_),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_1 _17808_ (.A0(net1827),
    .A1(_03890_),
    .S(_03915_),
    .X(_03917_));
 sky130_fd_sc_hd__clkbuf_1 _17809_ (.A(_03917_),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_1 _17810_ (.A0(\cur_mb_mem[206][2] ),
    .A1(_03892_),
    .S(_03915_),
    .X(_03918_));
 sky130_fd_sc_hd__clkbuf_1 _17811_ (.A(_03918_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _17812_ (.A0(\cur_mb_mem[206][3] ),
    .A1(_03894_),
    .S(_03915_),
    .X(_03919_));
 sky130_fd_sc_hd__clkbuf_1 _17813_ (.A(_03919_),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _17814_ (.A0(net1728),
    .A1(_03896_),
    .S(_03915_),
    .X(_03920_));
 sky130_fd_sc_hd__clkbuf_1 _17815_ (.A(_03920_),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_1 _17816_ (.A0(net1813),
    .A1(_03898_),
    .S(_03915_),
    .X(_03921_));
 sky130_fd_sc_hd__clkbuf_1 _17817_ (.A(_03921_),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _17818_ (.A0(\cur_mb_mem[206][6] ),
    .A1(_03900_),
    .S(_03915_),
    .X(_03922_));
 sky130_fd_sc_hd__clkbuf_1 _17819_ (.A(_03922_),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _17820_ (.A0(\cur_mb_mem[206][7] ),
    .A1(_03902_),
    .S(_03915_),
    .X(_03923_));
 sky130_fd_sc_hd__clkbuf_1 _17821_ (.A(_03923_),
    .X(_01806_));
 sky130_fd_sc_hd__and3_1 _17822_ (.A(_02406_),
    .B(_06094_),
    .C(_03826_),
    .X(_03924_));
 sky130_fd_sc_hd__clkbuf_8 _17823_ (.A(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__mux2_1 _17824_ (.A0(\cur_mb_mem[207][0] ),
    .A1(_03886_),
    .S(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__clkbuf_1 _17825_ (.A(_03926_),
    .X(_01807_));
 sky130_fd_sc_hd__mux2_1 _17826_ (.A0(\cur_mb_mem[207][1] ),
    .A1(_03890_),
    .S(_03925_),
    .X(_03927_));
 sky130_fd_sc_hd__clkbuf_1 _17827_ (.A(_03927_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _17828_ (.A0(net1868),
    .A1(_03892_),
    .S(_03925_),
    .X(_03928_));
 sky130_fd_sc_hd__clkbuf_1 _17829_ (.A(_03928_),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_1 _17830_ (.A0(\cur_mb_mem[207][3] ),
    .A1(_03894_),
    .S(_03925_),
    .X(_03929_));
 sky130_fd_sc_hd__clkbuf_1 _17831_ (.A(_03929_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _17832_ (.A0(\cur_mb_mem[207][4] ),
    .A1(_03896_),
    .S(_03925_),
    .X(_03930_));
 sky130_fd_sc_hd__clkbuf_1 _17833_ (.A(_03930_),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _17834_ (.A0(\cur_mb_mem[207][5] ),
    .A1(_03898_),
    .S(_03925_),
    .X(_03931_));
 sky130_fd_sc_hd__clkbuf_1 _17835_ (.A(_03931_),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _17836_ (.A0(\cur_mb_mem[207][6] ),
    .A1(_03900_),
    .S(_03925_),
    .X(_03932_));
 sky130_fd_sc_hd__clkbuf_1 _17837_ (.A(_03932_),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _17838_ (.A0(\cur_mb_mem[207][7] ),
    .A1(_03902_),
    .S(_03925_),
    .X(_03933_));
 sky130_fd_sc_hd__clkbuf_1 _17839_ (.A(_03933_),
    .X(_01814_));
 sky130_fd_sc_hd__clkbuf_4 _17840_ (.A(_06106_),
    .X(_03934_));
 sky130_fd_sc_hd__nand2_8 _17841_ (.A(_03934_),
    .B(_08882_),
    .Y(_03935_));
 sky130_fd_sc_hd__mux2_1 _17842_ (.A0(_03674_),
    .A1(net1330),
    .S(_03935_),
    .X(_03936_));
 sky130_fd_sc_hd__clkbuf_1 _17843_ (.A(_03936_),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _17844_ (.A0(_03677_),
    .A1(net750),
    .S(_03935_),
    .X(_03937_));
 sky130_fd_sc_hd__clkbuf_1 _17845_ (.A(_03937_),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _17846_ (.A0(_03679_),
    .A1(net512),
    .S(_03935_),
    .X(_03938_));
 sky130_fd_sc_hd__clkbuf_1 _17847_ (.A(_03938_),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _17848_ (.A0(_03681_),
    .A1(net1053),
    .S(_03935_),
    .X(_03939_));
 sky130_fd_sc_hd__clkbuf_1 _17849_ (.A(_03939_),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _17850_ (.A0(_03683_),
    .A1(net1032),
    .S(_03935_),
    .X(_03940_));
 sky130_fd_sc_hd__clkbuf_1 _17851_ (.A(_03940_),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _17852_ (.A0(_03685_),
    .A1(net1593),
    .S(_03935_),
    .X(_03941_));
 sky130_fd_sc_hd__clkbuf_1 _17853_ (.A(_03941_),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _17854_ (.A0(_03687_),
    .A1(net1321),
    .S(_03935_),
    .X(_03942_));
 sky130_fd_sc_hd__clkbuf_1 _17855_ (.A(_03942_),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_1 _17856_ (.A0(_03689_),
    .A1(net1028),
    .S(_03935_),
    .X(_03943_));
 sky130_fd_sc_hd__clkbuf_1 _17857_ (.A(_03943_),
    .X(_01822_));
 sky130_fd_sc_hd__nand2_4 _17858_ (.A(_06271_),
    .B(_03605_),
    .Y(_03944_));
 sky130_fd_sc_hd__mux2_1 _17859_ (.A0(_03674_),
    .A1(net1088),
    .S(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__clkbuf_1 _17860_ (.A(_03945_),
    .X(_01823_));
 sky130_fd_sc_hd__mux2_1 _17861_ (.A0(_03677_),
    .A1(net1808),
    .S(_03944_),
    .X(_03946_));
 sky130_fd_sc_hd__clkbuf_1 _17862_ (.A(_03946_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _17863_ (.A0(_03679_),
    .A1(net1176),
    .S(_03944_),
    .X(_03947_));
 sky130_fd_sc_hd__clkbuf_1 _17864_ (.A(_03947_),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _17865_ (.A0(_03681_),
    .A1(net602),
    .S(_03944_),
    .X(_03948_));
 sky130_fd_sc_hd__clkbuf_1 _17866_ (.A(_03948_),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_1 _17867_ (.A0(_03683_),
    .A1(net1935),
    .S(_03944_),
    .X(_03949_));
 sky130_fd_sc_hd__clkbuf_1 _17868_ (.A(_03949_),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _17869_ (.A0(_03685_),
    .A1(net1810),
    .S(_03944_),
    .X(_03950_));
 sky130_fd_sc_hd__clkbuf_1 _17870_ (.A(_03950_),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_1 _17871_ (.A0(_03687_),
    .A1(\cur_mb_mem[209][6] ),
    .S(_03944_),
    .X(_03951_));
 sky130_fd_sc_hd__clkbuf_1 _17872_ (.A(_03951_),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _17873_ (.A0(_03689_),
    .A1(net1850),
    .S(_03944_),
    .X(_03952_));
 sky130_fd_sc_hd__clkbuf_1 _17874_ (.A(_03952_),
    .X(_01830_));
 sky130_fd_sc_hd__nand2_8 _17875_ (.A(_06342_),
    .B(_03605_),
    .Y(_03953_));
 sky130_fd_sc_hd__mux2_1 _17876_ (.A0(_03674_),
    .A1(net635),
    .S(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__clkbuf_1 _17877_ (.A(_03954_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _17878_ (.A0(_03677_),
    .A1(net1205),
    .S(_03953_),
    .X(_03955_));
 sky130_fd_sc_hd__clkbuf_1 _17879_ (.A(_03955_),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _17880_ (.A0(_03679_),
    .A1(net1143),
    .S(_03953_),
    .X(_03956_));
 sky130_fd_sc_hd__clkbuf_1 _17881_ (.A(_03956_),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _17882_ (.A0(_03681_),
    .A1(net569),
    .S(_03953_),
    .X(_03957_));
 sky130_fd_sc_hd__clkbuf_1 _17883_ (.A(_03957_),
    .X(_01834_));
 sky130_fd_sc_hd__mux2_1 _17884_ (.A0(_03683_),
    .A1(net790),
    .S(_03953_),
    .X(_03958_));
 sky130_fd_sc_hd__clkbuf_1 _17885_ (.A(_03958_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _17886_ (.A0(_03685_),
    .A1(net668),
    .S(_03953_),
    .X(_03959_));
 sky130_fd_sc_hd__clkbuf_1 _17887_ (.A(_03959_),
    .X(_01836_));
 sky130_fd_sc_hd__mux2_1 _17888_ (.A0(_03687_),
    .A1(net1184),
    .S(_03953_),
    .X(_03960_));
 sky130_fd_sc_hd__clkbuf_1 _17889_ (.A(_03960_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _17890_ (.A0(_03689_),
    .A1(net1248),
    .S(_03953_),
    .X(_03961_));
 sky130_fd_sc_hd__clkbuf_1 _17891_ (.A(_03961_),
    .X(_01838_));
 sky130_fd_sc_hd__and3_1 _17892_ (.A(_02266_),
    .B(_03934_),
    .C(_03826_),
    .X(_03962_));
 sky130_fd_sc_hd__buf_4 _17893_ (.A(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__mux2_1 _17894_ (.A0(\cur_mb_mem[211][0] ),
    .A1(_03886_),
    .S(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__clkbuf_1 _17895_ (.A(_03964_),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_1 _17896_ (.A0(\cur_mb_mem[211][1] ),
    .A1(_03890_),
    .S(_03963_),
    .X(_03965_));
 sky130_fd_sc_hd__clkbuf_1 _17897_ (.A(_03965_),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _17898_ (.A0(\cur_mb_mem[211][2] ),
    .A1(_03892_),
    .S(_03963_),
    .X(_03966_));
 sky130_fd_sc_hd__clkbuf_1 _17899_ (.A(_03966_),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _17900_ (.A0(\cur_mb_mem[211][3] ),
    .A1(_03894_),
    .S(_03963_),
    .X(_03967_));
 sky130_fd_sc_hd__clkbuf_1 _17901_ (.A(_03967_),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _17902_ (.A0(net1105),
    .A1(_03896_),
    .S(_03963_),
    .X(_03968_));
 sky130_fd_sc_hd__clkbuf_1 _17903_ (.A(_03968_),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _17904_ (.A0(net1522),
    .A1(_03898_),
    .S(_03963_),
    .X(_03969_));
 sky130_fd_sc_hd__clkbuf_1 _17905_ (.A(_03969_),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _17906_ (.A0(\cur_mb_mem[211][6] ),
    .A1(_03900_),
    .S(_03963_),
    .X(_03970_));
 sky130_fd_sc_hd__clkbuf_1 _17907_ (.A(_03970_),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _17908_ (.A0(\cur_mb_mem[211][7] ),
    .A1(_03902_),
    .S(_03963_),
    .X(_03971_));
 sky130_fd_sc_hd__clkbuf_1 _17909_ (.A(_03971_),
    .X(_01846_));
 sky130_fd_sc_hd__nand2_8 _17910_ (.A(_06135_),
    .B(_03605_),
    .Y(_03972_));
 sky130_fd_sc_hd__mux2_1 _17911_ (.A0(_03674_),
    .A1(net1917),
    .S(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__clkbuf_1 _17912_ (.A(_03973_),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _17913_ (.A0(_03677_),
    .A1(net911),
    .S(_03972_),
    .X(_03974_));
 sky130_fd_sc_hd__clkbuf_1 _17914_ (.A(_03974_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _17915_ (.A0(_03679_),
    .A1(net907),
    .S(_03972_),
    .X(_03975_));
 sky130_fd_sc_hd__clkbuf_1 _17916_ (.A(_03975_),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _17917_ (.A0(_03681_),
    .A1(net559),
    .S(_03972_),
    .X(_03976_));
 sky130_fd_sc_hd__clkbuf_1 _17918_ (.A(_03976_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _17919_ (.A0(_03683_),
    .A1(net1122),
    .S(_03972_),
    .X(_03977_));
 sky130_fd_sc_hd__clkbuf_1 _17920_ (.A(_03977_),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _17921_ (.A0(_03685_),
    .A1(net983),
    .S(_03972_),
    .X(_03978_));
 sky130_fd_sc_hd__clkbuf_1 _17922_ (.A(_03978_),
    .X(_01852_));
 sky130_fd_sc_hd__mux2_1 _17923_ (.A0(_03687_),
    .A1(\cur_mb_mem[212][6] ),
    .S(_03972_),
    .X(_03979_));
 sky130_fd_sc_hd__clkbuf_1 _17924_ (.A(_03979_),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _17925_ (.A0(_03689_),
    .A1(net1312),
    .S(_03972_),
    .X(_03980_));
 sky130_fd_sc_hd__clkbuf_1 _17926_ (.A(_03980_),
    .X(_01854_));
 sky130_fd_sc_hd__clkbuf_2 _17927_ (.A(_08880_),
    .X(_03981_));
 sky130_fd_sc_hd__and3_1 _17928_ (.A(_03934_),
    .B(_02286_),
    .C(_03981_),
    .X(_03982_));
 sky130_fd_sc_hd__buf_4 _17929_ (.A(_03982_),
    .X(_03983_));
 sky130_fd_sc_hd__mux2_1 _17930_ (.A0(\cur_mb_mem[213][0] ),
    .A1(_03886_),
    .S(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__clkbuf_1 _17931_ (.A(_03984_),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _17932_ (.A0(\cur_mb_mem[213][1] ),
    .A1(_03890_),
    .S(_03983_),
    .X(_03985_));
 sky130_fd_sc_hd__clkbuf_1 _17933_ (.A(_03985_),
    .X(_01856_));
 sky130_fd_sc_hd__mux2_1 _17934_ (.A0(\cur_mb_mem[213][2] ),
    .A1(_03892_),
    .S(_03983_),
    .X(_03986_));
 sky130_fd_sc_hd__clkbuf_1 _17935_ (.A(_03986_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _17936_ (.A0(net1660),
    .A1(_03894_),
    .S(_03983_),
    .X(_03987_));
 sky130_fd_sc_hd__clkbuf_1 _17937_ (.A(_03987_),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _17938_ (.A0(net1955),
    .A1(_03896_),
    .S(_03983_),
    .X(_03988_));
 sky130_fd_sc_hd__clkbuf_1 _17939_ (.A(_03988_),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_1 _17940_ (.A0(net1956),
    .A1(_03898_),
    .S(_03983_),
    .X(_03989_));
 sky130_fd_sc_hd__clkbuf_1 _17941_ (.A(_03989_),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_1 _17942_ (.A0(\cur_mb_mem[213][6] ),
    .A1(_03900_),
    .S(_03983_),
    .X(_03990_));
 sky130_fd_sc_hd__clkbuf_1 _17943_ (.A(_03990_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _17944_ (.A0(net1874),
    .A1(_03902_),
    .S(_03983_),
    .X(_03991_));
 sky130_fd_sc_hd__clkbuf_1 _17945_ (.A(_03991_),
    .X(_01862_));
 sky130_fd_sc_hd__and3_1 _17946_ (.A(_02297_),
    .B(_03934_),
    .C(_03981_),
    .X(_03992_));
 sky130_fd_sc_hd__buf_4 _17947_ (.A(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__mux2_1 _17948_ (.A0(net1889),
    .A1(_03886_),
    .S(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__clkbuf_1 _17949_ (.A(_03994_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _17950_ (.A0(\cur_mb_mem[214][1] ),
    .A1(_03890_),
    .S(_03993_),
    .X(_03995_));
 sky130_fd_sc_hd__clkbuf_1 _17951_ (.A(_03995_),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _17952_ (.A0(net1859),
    .A1(_03892_),
    .S(_03993_),
    .X(_03996_));
 sky130_fd_sc_hd__clkbuf_1 _17953_ (.A(_03996_),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _17954_ (.A0(net1697),
    .A1(_03894_),
    .S(_03993_),
    .X(_03997_));
 sky130_fd_sc_hd__clkbuf_1 _17955_ (.A(_03997_),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _17956_ (.A0(net1951),
    .A1(_03896_),
    .S(_03993_),
    .X(_03998_));
 sky130_fd_sc_hd__clkbuf_1 _17957_ (.A(_03998_),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _17958_ (.A0(net1965),
    .A1(_03898_),
    .S(_03993_),
    .X(_03999_));
 sky130_fd_sc_hd__clkbuf_1 _17959_ (.A(_03999_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _17960_ (.A0(\cur_mb_mem[214][6] ),
    .A1(_03900_),
    .S(_03993_),
    .X(_04000_));
 sky130_fd_sc_hd__clkbuf_1 _17961_ (.A(_04000_),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _17962_ (.A0(\cur_mb_mem[214][7] ),
    .A1(_03902_),
    .S(_03993_),
    .X(_04001_));
 sky130_fd_sc_hd__clkbuf_1 _17963_ (.A(_04001_),
    .X(_01870_));
 sky130_fd_sc_hd__and3_1 _17964_ (.A(_03934_),
    .B(_06103_),
    .C(_03981_),
    .X(_04002_));
 sky130_fd_sc_hd__buf_4 _17965_ (.A(_04002_),
    .X(_04003_));
 sky130_fd_sc_hd__mux2_1 _17966_ (.A0(\cur_mb_mem[215][0] ),
    .A1(_03886_),
    .S(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__clkbuf_1 _17967_ (.A(_04004_),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _17968_ (.A0(\cur_mb_mem[215][1] ),
    .A1(_03890_),
    .S(_04003_),
    .X(_04005_));
 sky130_fd_sc_hd__clkbuf_1 _17969_ (.A(_04005_),
    .X(_01872_));
 sky130_fd_sc_hd__mux2_1 _17970_ (.A0(\cur_mb_mem[215][2] ),
    .A1(_03892_),
    .S(_04003_),
    .X(_04006_));
 sky130_fd_sc_hd__clkbuf_1 _17971_ (.A(_04006_),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _17972_ (.A0(\cur_mb_mem[215][3] ),
    .A1(_03894_),
    .S(_04003_),
    .X(_04007_));
 sky130_fd_sc_hd__clkbuf_1 _17973_ (.A(_04007_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _17974_ (.A0(\cur_mb_mem[215][4] ),
    .A1(_03896_),
    .S(_04003_),
    .X(_04008_));
 sky130_fd_sc_hd__clkbuf_1 _17975_ (.A(_04008_),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _17976_ (.A0(\cur_mb_mem[215][5] ),
    .A1(_03898_),
    .S(_04003_),
    .X(_04009_));
 sky130_fd_sc_hd__clkbuf_1 _17977_ (.A(_04009_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _17978_ (.A0(\cur_mb_mem[215][6] ),
    .A1(_03900_),
    .S(_04003_),
    .X(_04010_));
 sky130_fd_sc_hd__clkbuf_1 _17979_ (.A(_04010_),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _17980_ (.A0(net1990),
    .A1(_03902_),
    .S(_04003_),
    .X(_04011_));
 sky130_fd_sc_hd__clkbuf_1 _17981_ (.A(_04011_),
    .X(_01878_));
 sky130_fd_sc_hd__buf_2 _17982_ (.A(net97),
    .X(_04012_));
 sky130_fd_sc_hd__nand2_4 _17983_ (.A(_06317_),
    .B(_08979_),
    .Y(_04013_));
 sky130_fd_sc_hd__mux2_1 _17984_ (.A0(_04012_),
    .A1(net1632),
    .S(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__clkbuf_1 _17985_ (.A(_04014_),
    .X(_01879_));
 sky130_fd_sc_hd__clkbuf_4 _17986_ (.A(net98),
    .X(_04015_));
 sky130_fd_sc_hd__mux2_1 _17987_ (.A0(_04015_),
    .A1(\cur_mb_mem[216][1] ),
    .S(_04013_),
    .X(_04016_));
 sky130_fd_sc_hd__clkbuf_1 _17988_ (.A(_04016_),
    .X(_01880_));
 sky130_fd_sc_hd__clkbuf_4 _17989_ (.A(net99),
    .X(_04017_));
 sky130_fd_sc_hd__mux2_1 _17990_ (.A0(_04017_),
    .A1(net1561),
    .S(_04013_),
    .X(_04018_));
 sky130_fd_sc_hd__clkbuf_1 _17991_ (.A(_04018_),
    .X(_01881_));
 sky130_fd_sc_hd__clkbuf_4 _17992_ (.A(net100),
    .X(_04019_));
 sky130_fd_sc_hd__mux2_1 _17993_ (.A0(_04019_),
    .A1(net1678),
    .S(_04013_),
    .X(_04020_));
 sky130_fd_sc_hd__clkbuf_1 _17994_ (.A(_04020_),
    .X(_01882_));
 sky130_fd_sc_hd__buf_4 _17995_ (.A(net101),
    .X(_04021_));
 sky130_fd_sc_hd__mux2_1 _17996_ (.A0(_04021_),
    .A1(\cur_mb_mem[216][4] ),
    .S(_04013_),
    .X(_04022_));
 sky130_fd_sc_hd__clkbuf_1 _17997_ (.A(_04022_),
    .X(_01883_));
 sky130_fd_sc_hd__clkbuf_4 _17998_ (.A(net102),
    .X(_04023_));
 sky130_fd_sc_hd__mux2_1 _17999_ (.A0(_04023_),
    .A1(\cur_mb_mem[216][5] ),
    .S(_04013_),
    .X(_04024_));
 sky130_fd_sc_hd__clkbuf_1 _18000_ (.A(_04024_),
    .X(_01884_));
 sky130_fd_sc_hd__clkbuf_4 _18001_ (.A(net103),
    .X(_04025_));
 sky130_fd_sc_hd__mux2_1 _18002_ (.A0(_04025_),
    .A1(\cur_mb_mem[216][6] ),
    .S(_04013_),
    .X(_04026_));
 sky130_fd_sc_hd__clkbuf_1 _18003_ (.A(_04026_),
    .X(_01885_));
 sky130_fd_sc_hd__buf_4 _18004_ (.A(net104),
    .X(_04027_));
 sky130_fd_sc_hd__mux2_1 _18005_ (.A0(_04027_),
    .A1(\cur_mb_mem[216][7] ),
    .S(_04013_),
    .X(_04028_));
 sky130_fd_sc_hd__clkbuf_1 _18006_ (.A(_04028_),
    .X(_01886_));
 sky130_fd_sc_hd__and3_1 _18007_ (.A(_08978_),
    .B(_03934_),
    .C(_03981_),
    .X(_04029_));
 sky130_fd_sc_hd__buf_4 _18008_ (.A(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__mux2_1 _18009_ (.A0(\cur_mb_mem[217][0] ),
    .A1(_03886_),
    .S(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__clkbuf_1 _18010_ (.A(_04031_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _18011_ (.A0(\cur_mb_mem[217][1] ),
    .A1(_03890_),
    .S(_04030_),
    .X(_04032_));
 sky130_fd_sc_hd__clkbuf_1 _18012_ (.A(_04032_),
    .X(_01888_));
 sky130_fd_sc_hd__mux2_1 _18013_ (.A0(net1901),
    .A1(_03892_),
    .S(_04030_),
    .X(_04033_));
 sky130_fd_sc_hd__clkbuf_1 _18014_ (.A(_04033_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _18015_ (.A0(net1119),
    .A1(_03894_),
    .S(_04030_),
    .X(_04034_));
 sky130_fd_sc_hd__clkbuf_1 _18016_ (.A(_04034_),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_1 _18017_ (.A0(net914),
    .A1(_03896_),
    .S(_04030_),
    .X(_04035_));
 sky130_fd_sc_hd__clkbuf_1 _18018_ (.A(_04035_),
    .X(_01891_));
 sky130_fd_sc_hd__mux2_1 _18019_ (.A0(net1364),
    .A1(_03898_),
    .S(_04030_),
    .X(_04036_));
 sky130_fd_sc_hd__clkbuf_1 _18020_ (.A(_04036_),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _18021_ (.A0(\cur_mb_mem[217][6] ),
    .A1(_03900_),
    .S(_04030_),
    .X(_04037_));
 sky130_fd_sc_hd__clkbuf_1 _18022_ (.A(_04037_),
    .X(_01893_));
 sky130_fd_sc_hd__mux2_1 _18023_ (.A0(\cur_mb_mem[217][7] ),
    .A1(_03902_),
    .S(_04030_),
    .X(_04038_));
 sky130_fd_sc_hd__clkbuf_1 _18024_ (.A(_04038_),
    .X(_01894_));
 sky130_fd_sc_hd__and3_1 _18025_ (.A(_02353_),
    .B(_03934_),
    .C(_03981_),
    .X(_04039_));
 sky130_fd_sc_hd__buf_4 _18026_ (.A(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__mux2_1 _18027_ (.A0(\cur_mb_mem[218][0] ),
    .A1(_03886_),
    .S(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__clkbuf_1 _18028_ (.A(_04041_),
    .X(_01895_));
 sky130_fd_sc_hd__mux2_1 _18029_ (.A0(\cur_mb_mem[218][1] ),
    .A1(_03890_),
    .S(_04040_),
    .X(_04042_));
 sky130_fd_sc_hd__clkbuf_1 _18030_ (.A(_04042_),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _18031_ (.A0(\cur_mb_mem[218][2] ),
    .A1(_03892_),
    .S(_04040_),
    .X(_04043_));
 sky130_fd_sc_hd__clkbuf_1 _18032_ (.A(_04043_),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _18033_ (.A0(net1699),
    .A1(_03894_),
    .S(_04040_),
    .X(_04044_));
 sky130_fd_sc_hd__clkbuf_1 _18034_ (.A(_04044_),
    .X(_01898_));
 sky130_fd_sc_hd__mux2_1 _18035_ (.A0(net1939),
    .A1(_03896_),
    .S(_04040_),
    .X(_04045_));
 sky130_fd_sc_hd__clkbuf_1 _18036_ (.A(_04045_),
    .X(_01899_));
 sky130_fd_sc_hd__mux2_1 _18037_ (.A0(net1970),
    .A1(_03898_),
    .S(_04040_),
    .X(_04046_));
 sky130_fd_sc_hd__clkbuf_1 _18038_ (.A(_04046_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_1 _18039_ (.A0(\cur_mb_mem[218][6] ),
    .A1(_03900_),
    .S(_04040_),
    .X(_04047_));
 sky130_fd_sc_hd__clkbuf_1 _18040_ (.A(_04047_),
    .X(_01901_));
 sky130_fd_sc_hd__mux2_1 _18041_ (.A0(\cur_mb_mem[218][7] ),
    .A1(_03902_),
    .S(_04040_),
    .X(_04048_));
 sky130_fd_sc_hd__clkbuf_1 _18042_ (.A(_04048_),
    .X(_01902_));
 sky130_fd_sc_hd__clkbuf_8 _18043_ (.A(_08530_),
    .X(_04049_));
 sky130_fd_sc_hd__and3_1 _18044_ (.A(_02526_),
    .B(_03934_),
    .C(_03981_),
    .X(_04050_));
 sky130_fd_sc_hd__clkbuf_8 _18045_ (.A(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__mux2_1 _18046_ (.A0(net1866),
    .A1(_04049_),
    .S(_04051_),
    .X(_04052_));
 sky130_fd_sc_hd__clkbuf_1 _18047_ (.A(_04052_),
    .X(_01903_));
 sky130_fd_sc_hd__buf_4 _18048_ (.A(_08535_),
    .X(_04053_));
 sky130_fd_sc_hd__mux2_1 _18049_ (.A0(net1040),
    .A1(_04053_),
    .S(_04051_),
    .X(_04054_));
 sky130_fd_sc_hd__clkbuf_1 _18050_ (.A(_04054_),
    .X(_01904_));
 sky130_fd_sc_hd__clkbuf_8 _18051_ (.A(_08538_),
    .X(_04055_));
 sky130_fd_sc_hd__mux2_1 _18052_ (.A0(net1771),
    .A1(_04055_),
    .S(_04051_),
    .X(_04056_));
 sky130_fd_sc_hd__clkbuf_1 _18053_ (.A(_04056_),
    .X(_01905_));
 sky130_fd_sc_hd__clkbuf_8 _18054_ (.A(_08541_),
    .X(_04057_));
 sky130_fd_sc_hd__mux2_1 _18055_ (.A0(net1869),
    .A1(_04057_),
    .S(_04051_),
    .X(_04058_));
 sky130_fd_sc_hd__clkbuf_1 _18056_ (.A(_04058_),
    .X(_01906_));
 sky130_fd_sc_hd__clkbuf_8 _18057_ (.A(_08544_),
    .X(_04059_));
 sky130_fd_sc_hd__mux2_1 _18058_ (.A0(\cur_mb_mem[219][4] ),
    .A1(_04059_),
    .S(_04051_),
    .X(_04060_));
 sky130_fd_sc_hd__clkbuf_1 _18059_ (.A(_04060_),
    .X(_01907_));
 sky130_fd_sc_hd__clkbuf_8 _18060_ (.A(_08547_),
    .X(_04061_));
 sky130_fd_sc_hd__mux2_1 _18061_ (.A0(net1709),
    .A1(_04061_),
    .S(_04051_),
    .X(_04062_));
 sky130_fd_sc_hd__clkbuf_1 _18062_ (.A(_04062_),
    .X(_01908_));
 sky130_fd_sc_hd__clkbuf_4 _18063_ (.A(_08550_),
    .X(_04063_));
 sky130_fd_sc_hd__mux2_1 _18064_ (.A0(\cur_mb_mem[219][6] ),
    .A1(_04063_),
    .S(_04051_),
    .X(_04064_));
 sky130_fd_sc_hd__clkbuf_1 _18065_ (.A(_04064_),
    .X(_01909_));
 sky130_fd_sc_hd__clkbuf_4 _18066_ (.A(_08553_),
    .X(_04065_));
 sky130_fd_sc_hd__mux2_1 _18067_ (.A0(\cur_mb_mem[219][7] ),
    .A1(_04065_),
    .S(_04051_),
    .X(_04066_));
 sky130_fd_sc_hd__clkbuf_1 _18068_ (.A(_04066_),
    .X(_01910_));
 sky130_fd_sc_hd__and3_1 _18069_ (.A(_02374_),
    .B(_03934_),
    .C(_03981_),
    .X(_04067_));
 sky130_fd_sc_hd__buf_4 _18070_ (.A(_04067_),
    .X(_04068_));
 sky130_fd_sc_hd__mux2_1 _18071_ (.A0(net641),
    .A1(_04049_),
    .S(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__clkbuf_1 _18072_ (.A(_04069_),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _18073_ (.A0(net744),
    .A1(_04053_),
    .S(_04068_),
    .X(_04070_));
 sky130_fd_sc_hd__clkbuf_1 _18074_ (.A(_04070_),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _18075_ (.A0(net832),
    .A1(_04055_),
    .S(_04068_),
    .X(_04071_));
 sky130_fd_sc_hd__clkbuf_1 _18076_ (.A(_04071_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _18077_ (.A0(net1552),
    .A1(_04057_),
    .S(_04068_),
    .X(_04072_));
 sky130_fd_sc_hd__clkbuf_1 _18078_ (.A(_04072_),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_1 _18079_ (.A0(net703),
    .A1(_04059_),
    .S(_04068_),
    .X(_04073_));
 sky130_fd_sc_hd__clkbuf_1 _18080_ (.A(_04073_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _18081_ (.A0(net751),
    .A1(_04061_),
    .S(_04068_),
    .X(_04074_));
 sky130_fd_sc_hd__clkbuf_1 _18082_ (.A(_04074_),
    .X(_01916_));
 sky130_fd_sc_hd__mux2_1 _18083_ (.A0(\cur_mb_mem[220][6] ),
    .A1(_04063_),
    .S(_04068_),
    .X(_04075_));
 sky130_fd_sc_hd__clkbuf_1 _18084_ (.A(_04075_),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_1 _18085_ (.A0(net1436),
    .A1(_04065_),
    .S(_04068_),
    .X(_04076_));
 sky130_fd_sc_hd__clkbuf_1 _18086_ (.A(_04076_),
    .X(_01918_));
 sky130_fd_sc_hd__and3_1 _18087_ (.A(_09025_),
    .B(_06106_),
    .C(_03981_),
    .X(_04077_));
 sky130_fd_sc_hd__buf_4 _18088_ (.A(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__mux2_1 _18089_ (.A0(net1727),
    .A1(_04049_),
    .S(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__clkbuf_1 _18090_ (.A(_04079_),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _18091_ (.A0(\cur_mb_mem[221][1] ),
    .A1(_04053_),
    .S(_04078_),
    .X(_04080_));
 sky130_fd_sc_hd__clkbuf_1 _18092_ (.A(_04080_),
    .X(_01920_));
 sky130_fd_sc_hd__mux2_1 _18093_ (.A0(net1653),
    .A1(_04055_),
    .S(_04078_),
    .X(_04081_));
 sky130_fd_sc_hd__clkbuf_1 _18094_ (.A(_04081_),
    .X(_01921_));
 sky130_fd_sc_hd__mux2_1 _18095_ (.A0(net1745),
    .A1(_04057_),
    .S(_04078_),
    .X(_04082_));
 sky130_fd_sc_hd__clkbuf_1 _18096_ (.A(_04082_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_1 _18097_ (.A0(net1957),
    .A1(_04059_),
    .S(_04078_),
    .X(_04083_));
 sky130_fd_sc_hd__clkbuf_1 _18098_ (.A(_04083_),
    .X(_01923_));
 sky130_fd_sc_hd__mux2_1 _18099_ (.A0(net1941),
    .A1(_04061_),
    .S(_04078_),
    .X(_04084_));
 sky130_fd_sc_hd__clkbuf_1 _18100_ (.A(_04084_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _18101_ (.A0(net1108),
    .A1(_04063_),
    .S(_04078_),
    .X(_04085_));
 sky130_fd_sc_hd__clkbuf_1 _18102_ (.A(_04085_),
    .X(_01925_));
 sky130_fd_sc_hd__mux2_1 _18103_ (.A0(net804),
    .A1(_04065_),
    .S(_04078_),
    .X(_04086_));
 sky130_fd_sc_hd__clkbuf_1 _18104_ (.A(_04086_),
    .X(_01926_));
 sky130_fd_sc_hd__and3_1 _18105_ (.A(_03934_),
    .B(_06025_),
    .C(_03981_),
    .X(_04087_));
 sky130_fd_sc_hd__buf_4 _18106_ (.A(_04087_),
    .X(_04088_));
 sky130_fd_sc_hd__mux2_1 _18107_ (.A0(net1509),
    .A1(_04049_),
    .S(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__clkbuf_1 _18108_ (.A(_04089_),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _18109_ (.A0(net586),
    .A1(_04053_),
    .S(_04088_),
    .X(_04090_));
 sky130_fd_sc_hd__clkbuf_1 _18110_ (.A(_04090_),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _18111_ (.A0(net923),
    .A1(_04055_),
    .S(_04088_),
    .X(_04091_));
 sky130_fd_sc_hd__clkbuf_1 _18112_ (.A(_04091_),
    .X(_01929_));
 sky130_fd_sc_hd__mux2_1 _18113_ (.A0(net1127),
    .A1(_04057_),
    .S(_04088_),
    .X(_04092_));
 sky130_fd_sc_hd__clkbuf_1 _18114_ (.A(_04092_),
    .X(_01930_));
 sky130_fd_sc_hd__mux2_1 _18115_ (.A0(net1918),
    .A1(_04059_),
    .S(_04088_),
    .X(_04093_));
 sky130_fd_sc_hd__clkbuf_1 _18116_ (.A(_04093_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_1 _18117_ (.A0(net1924),
    .A1(_04061_),
    .S(_04088_),
    .X(_04094_));
 sky130_fd_sc_hd__clkbuf_1 _18118_ (.A(_04094_),
    .X(_01932_));
 sky130_fd_sc_hd__mux2_1 _18119_ (.A0(\cur_mb_mem[222][6] ),
    .A1(_04063_),
    .S(_04088_),
    .X(_04095_));
 sky130_fd_sc_hd__clkbuf_1 _18120_ (.A(_04095_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _18121_ (.A0(net795),
    .A1(_04065_),
    .S(_04088_),
    .X(_04096_));
 sky130_fd_sc_hd__clkbuf_1 _18122_ (.A(_04096_),
    .X(_01934_));
 sky130_fd_sc_hd__and3_1 _18123_ (.A(_02406_),
    .B(_06106_),
    .C(_03981_),
    .X(_04097_));
 sky130_fd_sc_hd__buf_4 _18124_ (.A(_04097_),
    .X(_04098_));
 sky130_fd_sc_hd__mux2_1 _18125_ (.A0(\cur_mb_mem[223][0] ),
    .A1(_04049_),
    .S(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__clkbuf_1 _18126_ (.A(_04099_),
    .X(_01935_));
 sky130_fd_sc_hd__mux2_1 _18127_ (.A0(\cur_mb_mem[223][1] ),
    .A1(_04053_),
    .S(_04098_),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_1 _18128_ (.A(_04100_),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_1 _18129_ (.A0(\cur_mb_mem[223][2] ),
    .A1(_04055_),
    .S(_04098_),
    .X(_04101_));
 sky130_fd_sc_hd__clkbuf_1 _18130_ (.A(_04101_),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _18131_ (.A0(\cur_mb_mem[223][3] ),
    .A1(_04057_),
    .S(_04098_),
    .X(_04102_));
 sky130_fd_sc_hd__clkbuf_1 _18132_ (.A(_04102_),
    .X(_01938_));
 sky130_fd_sc_hd__mux2_1 _18133_ (.A0(\cur_mb_mem[223][4] ),
    .A1(_04059_),
    .S(_04098_),
    .X(_04103_));
 sky130_fd_sc_hd__clkbuf_1 _18134_ (.A(_04103_),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_1 _18135_ (.A0(\cur_mb_mem[223][5] ),
    .A1(_04061_),
    .S(_04098_),
    .X(_04104_));
 sky130_fd_sc_hd__clkbuf_1 _18136_ (.A(_04104_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_1 _18137_ (.A0(\cur_mb_mem[223][6] ),
    .A1(_04063_),
    .S(_04098_),
    .X(_04105_));
 sky130_fd_sc_hd__clkbuf_1 _18138_ (.A(_04105_),
    .X(_01941_));
 sky130_fd_sc_hd__mux2_1 _18139_ (.A0(\cur_mb_mem[223][7] ),
    .A1(_04065_),
    .S(_04098_),
    .X(_04106_));
 sky130_fd_sc_hd__clkbuf_1 _18140_ (.A(_04106_),
    .X(_01942_));
 sky130_fd_sc_hd__buf_4 _18141_ (.A(_06067_),
    .X(_04107_));
 sky130_fd_sc_hd__nand2_8 _18142_ (.A(_04107_),
    .B(_08882_),
    .Y(_04108_));
 sky130_fd_sc_hd__mux2_1 _18143_ (.A0(_04012_),
    .A1(net952),
    .S(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__clkbuf_1 _18144_ (.A(_04109_),
    .X(_01943_));
 sky130_fd_sc_hd__mux2_1 _18145_ (.A0(_04015_),
    .A1(\cur_mb_mem[224][1] ),
    .S(_04108_),
    .X(_04110_));
 sky130_fd_sc_hd__clkbuf_1 _18146_ (.A(_04110_),
    .X(_01944_));
 sky130_fd_sc_hd__mux2_1 _18147_ (.A0(_04017_),
    .A1(net1988),
    .S(_04108_),
    .X(_04111_));
 sky130_fd_sc_hd__clkbuf_1 _18148_ (.A(_04111_),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _18149_ (.A0(_04019_),
    .A1(net1915),
    .S(_04108_),
    .X(_04112_));
 sky130_fd_sc_hd__clkbuf_1 _18150_ (.A(_04112_),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _18151_ (.A0(_04021_),
    .A1(net1604),
    .S(_04108_),
    .X(_04113_));
 sky130_fd_sc_hd__clkbuf_1 _18152_ (.A(_04113_),
    .X(_01947_));
 sky130_fd_sc_hd__mux2_1 _18153_ (.A0(_04023_),
    .A1(net1562),
    .S(_04108_),
    .X(_04114_));
 sky130_fd_sc_hd__clkbuf_1 _18154_ (.A(_04114_),
    .X(_01948_));
 sky130_fd_sc_hd__mux2_1 _18155_ (.A0(_04025_),
    .A1(\cur_mb_mem[224][6] ),
    .S(_04108_),
    .X(_04115_));
 sky130_fd_sc_hd__clkbuf_1 _18156_ (.A(_04115_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _18157_ (.A0(_04027_),
    .A1(net1574),
    .S(_04108_),
    .X(_04116_));
 sky130_fd_sc_hd__clkbuf_1 _18158_ (.A(_04116_),
    .X(_01950_));
 sky130_fd_sc_hd__nand2_4 _18159_ (.A(_05998_),
    .B(_08979_),
    .Y(_04117_));
 sky130_fd_sc_hd__mux2_1 _18160_ (.A0(_04012_),
    .A1(\cur_mb_mem[225][0] ),
    .S(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_1 _18161_ (.A(_04118_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _18162_ (.A0(_04015_),
    .A1(net1297),
    .S(_04117_),
    .X(_04119_));
 sky130_fd_sc_hd__clkbuf_1 _18163_ (.A(_04119_),
    .X(_01952_));
 sky130_fd_sc_hd__mux2_1 _18164_ (.A0(_04017_),
    .A1(\cur_mb_mem[225][2] ),
    .S(_04117_),
    .X(_04120_));
 sky130_fd_sc_hd__clkbuf_1 _18165_ (.A(_04120_),
    .X(_01953_));
 sky130_fd_sc_hd__mux2_1 _18166_ (.A0(_04019_),
    .A1(\cur_mb_mem[225][3] ),
    .S(_04117_),
    .X(_04121_));
 sky130_fd_sc_hd__clkbuf_1 _18167_ (.A(_04121_),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _18168_ (.A0(_04021_),
    .A1(net1486),
    .S(_04117_),
    .X(_04122_));
 sky130_fd_sc_hd__clkbuf_1 _18169_ (.A(_04122_),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _18170_ (.A0(_04023_),
    .A1(net1523),
    .S(_04117_),
    .X(_04123_));
 sky130_fd_sc_hd__clkbuf_1 _18171_ (.A(_04123_),
    .X(_01956_));
 sky130_fd_sc_hd__mux2_1 _18172_ (.A0(_04025_),
    .A1(\cur_mb_mem[225][6] ),
    .S(_04117_),
    .X(_04124_));
 sky130_fd_sc_hd__clkbuf_1 _18173_ (.A(_04124_),
    .X(_01957_));
 sky130_fd_sc_hd__mux2_1 _18174_ (.A0(_04027_),
    .A1(\cur_mb_mem[225][7] ),
    .S(_04117_),
    .X(_04125_));
 sky130_fd_sc_hd__clkbuf_1 _18175_ (.A(_04125_),
    .X(_01958_));
 sky130_fd_sc_hd__nand2_4 _18176_ (.A(_06256_),
    .B(_08979_),
    .Y(_04126_));
 sky130_fd_sc_hd__mux2_1 _18177_ (.A0(_04012_),
    .A1(net1251),
    .S(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__clkbuf_1 _18178_ (.A(_04127_),
    .X(_01959_));
 sky130_fd_sc_hd__mux2_1 _18179_ (.A0(_04015_),
    .A1(\cur_mb_mem[226][1] ),
    .S(_04126_),
    .X(_04128_));
 sky130_fd_sc_hd__clkbuf_1 _18180_ (.A(_04128_),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_1 _18181_ (.A0(_04017_),
    .A1(net1303),
    .S(_04126_),
    .X(_04129_));
 sky130_fd_sc_hd__clkbuf_1 _18182_ (.A(_04129_),
    .X(_01961_));
 sky130_fd_sc_hd__mux2_1 _18183_ (.A0(_04019_),
    .A1(net1346),
    .S(_04126_),
    .X(_04130_));
 sky130_fd_sc_hd__clkbuf_1 _18184_ (.A(_04130_),
    .X(_01962_));
 sky130_fd_sc_hd__mux2_1 _18185_ (.A0(_04021_),
    .A1(net1714),
    .S(_04126_),
    .X(_04131_));
 sky130_fd_sc_hd__clkbuf_1 _18186_ (.A(_04131_),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _18187_ (.A0(_04023_),
    .A1(net1763),
    .S(_04126_),
    .X(_04132_));
 sky130_fd_sc_hd__clkbuf_1 _18188_ (.A(_04132_),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _18189_ (.A0(_04025_),
    .A1(\cur_mb_mem[226][6] ),
    .S(_04126_),
    .X(_04133_));
 sky130_fd_sc_hd__clkbuf_1 _18190_ (.A(_04133_),
    .X(_01965_));
 sky130_fd_sc_hd__mux2_1 _18191_ (.A0(_04027_),
    .A1(\cur_mb_mem[226][7] ),
    .S(_04126_),
    .X(_04134_));
 sky130_fd_sc_hd__clkbuf_1 _18192_ (.A(_04134_),
    .X(_01966_));
 sky130_fd_sc_hd__buf_2 _18193_ (.A(_08880_),
    .X(_04135_));
 sky130_fd_sc_hd__and3_1 _18194_ (.A(_02266_),
    .B(_04107_),
    .C(_04135_),
    .X(_04136_));
 sky130_fd_sc_hd__buf_4 _18195_ (.A(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__mux2_1 _18196_ (.A0(\cur_mb_mem[227][0] ),
    .A1(_04049_),
    .S(_04137_),
    .X(_04138_));
 sky130_fd_sc_hd__clkbuf_1 _18197_ (.A(_04138_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _18198_ (.A0(net1919),
    .A1(_04053_),
    .S(_04137_),
    .X(_04139_));
 sky130_fd_sc_hd__clkbuf_1 _18199_ (.A(_04139_),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_1 _18200_ (.A0(\cur_mb_mem[227][2] ),
    .A1(_04055_),
    .S(_04137_),
    .X(_04140_));
 sky130_fd_sc_hd__clkbuf_1 _18201_ (.A(_04140_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _18202_ (.A0(net1543),
    .A1(_04057_),
    .S(_04137_),
    .X(_04141_));
 sky130_fd_sc_hd__clkbuf_1 _18203_ (.A(_04141_),
    .X(_01970_));
 sky130_fd_sc_hd__mux2_1 _18204_ (.A0(net1111),
    .A1(_04059_),
    .S(_04137_),
    .X(_04142_));
 sky130_fd_sc_hd__clkbuf_1 _18205_ (.A(_04142_),
    .X(_01971_));
 sky130_fd_sc_hd__mux2_1 _18206_ (.A0(net757),
    .A1(_04061_),
    .S(_04137_),
    .X(_04143_));
 sky130_fd_sc_hd__clkbuf_1 _18207_ (.A(_04143_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _18208_ (.A0(net1886),
    .A1(_04063_),
    .S(_04137_),
    .X(_04144_));
 sky130_fd_sc_hd__clkbuf_1 _18209_ (.A(_04144_),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _18210_ (.A0(net949),
    .A1(_04065_),
    .S(_04137_),
    .X(_04145_));
 sky130_fd_sc_hd__clkbuf_1 _18211_ (.A(_04145_),
    .X(_01974_));
 sky130_fd_sc_hd__nand3_4 _18212_ (.A(_06223_),
    .B(_04107_),
    .C(_08901_),
    .Y(_04146_));
 sky130_fd_sc_hd__mux2_1 _18213_ (.A0(_04012_),
    .A1(\cur_mb_mem[228][0] ),
    .S(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__clkbuf_1 _18214_ (.A(_04147_),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_1 _18215_ (.A0(_04015_),
    .A1(\cur_mb_mem[228][1] ),
    .S(_04146_),
    .X(_04148_));
 sky130_fd_sc_hd__clkbuf_1 _18216_ (.A(_04148_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_1 _18217_ (.A0(_04017_),
    .A1(net1837),
    .S(_04146_),
    .X(_04149_));
 sky130_fd_sc_hd__clkbuf_1 _18218_ (.A(_04149_),
    .X(_01977_));
 sky130_fd_sc_hd__mux2_1 _18219_ (.A0(_04019_),
    .A1(net1896),
    .S(_04146_),
    .X(_04150_));
 sky130_fd_sc_hd__clkbuf_1 _18220_ (.A(_04150_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _18221_ (.A0(_04021_),
    .A1(net1920),
    .S(_04146_),
    .X(_04151_));
 sky130_fd_sc_hd__clkbuf_1 _18222_ (.A(_04151_),
    .X(_01979_));
 sky130_fd_sc_hd__mux2_1 _18223_ (.A0(_04023_),
    .A1(net1856),
    .S(_04146_),
    .X(_04152_));
 sky130_fd_sc_hd__clkbuf_1 _18224_ (.A(_04152_),
    .X(_01980_));
 sky130_fd_sc_hd__mux2_1 _18225_ (.A0(_04025_),
    .A1(\cur_mb_mem[228][6] ),
    .S(_04146_),
    .X(_04153_));
 sky130_fd_sc_hd__clkbuf_1 _18226_ (.A(_04153_),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _18227_ (.A0(_04027_),
    .A1(net1357),
    .S(_04146_),
    .X(_04154_));
 sky130_fd_sc_hd__clkbuf_1 _18228_ (.A(_04154_),
    .X(_01982_));
 sky130_fd_sc_hd__and3_1 _18229_ (.A(_02286_),
    .B(_04107_),
    .C(_04135_),
    .X(_04155_));
 sky130_fd_sc_hd__clkbuf_4 _18230_ (.A(_04155_),
    .X(_04156_));
 sky130_fd_sc_hd__mux2_1 _18231_ (.A0(net817),
    .A1(_04049_),
    .S(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__clkbuf_1 _18232_ (.A(_04157_),
    .X(_01983_));
 sky130_fd_sc_hd__mux2_1 _18233_ (.A0(net682),
    .A1(_04053_),
    .S(_04156_),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_1 _18234_ (.A(_04158_),
    .X(_01984_));
 sky130_fd_sc_hd__mux2_1 _18235_ (.A0(net874),
    .A1(_04055_),
    .S(_04156_),
    .X(_04159_));
 sky130_fd_sc_hd__clkbuf_1 _18236_ (.A(_04159_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _18237_ (.A0(net828),
    .A1(_04057_),
    .S(_04156_),
    .X(_04160_));
 sky130_fd_sc_hd__clkbuf_1 _18238_ (.A(_04160_),
    .X(_01986_));
 sky130_fd_sc_hd__mux2_1 _18239_ (.A0(net526),
    .A1(_04059_),
    .S(_04156_),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_1 _18240_ (.A(_04161_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _18241_ (.A0(net1566),
    .A1(_04061_),
    .S(_04156_),
    .X(_04162_));
 sky130_fd_sc_hd__clkbuf_1 _18242_ (.A(_04162_),
    .X(_01988_));
 sky130_fd_sc_hd__mux2_1 _18243_ (.A0(\cur_mb_mem[229][6] ),
    .A1(_04063_),
    .S(_04156_),
    .X(_04163_));
 sky130_fd_sc_hd__clkbuf_1 _18244_ (.A(_04163_),
    .X(_01989_));
 sky130_fd_sc_hd__mux2_1 _18245_ (.A0(net333),
    .A1(_04065_),
    .S(_04156_),
    .X(_04164_));
 sky130_fd_sc_hd__clkbuf_1 _18246_ (.A(_04164_),
    .X(_01990_));
 sky130_fd_sc_hd__and3_1 _18247_ (.A(_02297_),
    .B(_04107_),
    .C(_04135_),
    .X(_04165_));
 sky130_fd_sc_hd__buf_4 _18248_ (.A(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__mux2_1 _18249_ (.A0(net1659),
    .A1(_04049_),
    .S(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__clkbuf_1 _18250_ (.A(_04167_),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _18251_ (.A0(net1744),
    .A1(_04053_),
    .S(_04166_),
    .X(_04168_));
 sky130_fd_sc_hd__clkbuf_1 _18252_ (.A(_04168_),
    .X(_01992_));
 sky130_fd_sc_hd__mux2_1 _18253_ (.A0(net606),
    .A1(_04055_),
    .S(_04166_),
    .X(_04169_));
 sky130_fd_sc_hd__clkbuf_1 _18254_ (.A(_04169_),
    .X(_01993_));
 sky130_fd_sc_hd__mux2_1 _18255_ (.A0(net1927),
    .A1(_04057_),
    .S(_04166_),
    .X(_04170_));
 sky130_fd_sc_hd__clkbuf_1 _18256_ (.A(_04170_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_1 _18257_ (.A0(net615),
    .A1(_04059_),
    .S(_04166_),
    .X(_04171_));
 sky130_fd_sc_hd__clkbuf_1 _18258_ (.A(_04171_),
    .X(_01995_));
 sky130_fd_sc_hd__mux2_1 _18259_ (.A0(net865),
    .A1(_04061_),
    .S(_04166_),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _18260_ (.A(_04172_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _18261_ (.A0(net991),
    .A1(_04063_),
    .S(_04166_),
    .X(_04173_));
 sky130_fd_sc_hd__clkbuf_1 _18262_ (.A(_04173_),
    .X(_01997_));
 sky130_fd_sc_hd__mux2_1 _18263_ (.A0(net437),
    .A1(_04065_),
    .S(_04166_),
    .X(_04174_));
 sky130_fd_sc_hd__clkbuf_1 _18264_ (.A(_04174_),
    .X(_01998_));
 sky130_fd_sc_hd__and3_1 _18265_ (.A(_08839_),
    .B(_04107_),
    .C(_04135_),
    .X(_04175_));
 sky130_fd_sc_hd__buf_4 _18266_ (.A(_04175_),
    .X(_04176_));
 sky130_fd_sc_hd__mux2_1 _18267_ (.A0(\cur_mb_mem[231][0] ),
    .A1(_04049_),
    .S(_04176_),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_1 _18268_ (.A(_04177_),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _18269_ (.A0(net1770),
    .A1(_04053_),
    .S(_04176_),
    .X(_04178_));
 sky130_fd_sc_hd__clkbuf_1 _18270_ (.A(_04178_),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_1 _18271_ (.A0(\cur_mb_mem[231][2] ),
    .A1(_04055_),
    .S(_04176_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _18272_ (.A(_04179_),
    .X(_02001_));
 sky130_fd_sc_hd__mux2_1 _18273_ (.A0(\cur_mb_mem[231][3] ),
    .A1(_04057_),
    .S(_04176_),
    .X(_04180_));
 sky130_fd_sc_hd__clkbuf_1 _18274_ (.A(_04180_),
    .X(_02002_));
 sky130_fd_sc_hd__mux2_1 _18275_ (.A0(net1823),
    .A1(_04059_),
    .S(_04176_),
    .X(_04181_));
 sky130_fd_sc_hd__clkbuf_1 _18276_ (.A(_04181_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_1 _18277_ (.A0(net1296),
    .A1(_04061_),
    .S(_04176_),
    .X(_04182_));
 sky130_fd_sc_hd__clkbuf_1 _18278_ (.A(_04182_),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_1 _18279_ (.A0(\cur_mb_mem[231][6] ),
    .A1(_04063_),
    .S(_04176_),
    .X(_04183_));
 sky130_fd_sc_hd__clkbuf_1 _18280_ (.A(_04183_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _18281_ (.A0(\cur_mb_mem[231][7] ),
    .A1(_04065_),
    .S(_04176_),
    .X(_04184_));
 sky130_fd_sc_hd__clkbuf_1 _18282_ (.A(_04184_),
    .X(_02006_));
 sky130_fd_sc_hd__nand2_4 _18283_ (.A(_06463_),
    .B(_08979_),
    .Y(_04185_));
 sky130_fd_sc_hd__mux2_1 _18284_ (.A0(_04012_),
    .A1(net1982),
    .S(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__clkbuf_1 _18285_ (.A(_04186_),
    .X(_02007_));
 sky130_fd_sc_hd__mux2_1 _18286_ (.A0(_04015_),
    .A1(net1821),
    .S(_04185_),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_1 _18287_ (.A(_04187_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _18288_ (.A0(_04017_),
    .A1(net1739),
    .S(_04185_),
    .X(_04188_));
 sky130_fd_sc_hd__clkbuf_1 _18289_ (.A(_04188_),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _18290_ (.A0(_04019_),
    .A1(net1765),
    .S(_04185_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _18291_ (.A(_04189_),
    .X(_02010_));
 sky130_fd_sc_hd__mux2_1 _18292_ (.A0(_04021_),
    .A1(net1736),
    .S(_04185_),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_1 _18293_ (.A(_04190_),
    .X(_02011_));
 sky130_fd_sc_hd__mux2_1 _18294_ (.A0(_04023_),
    .A1(net1841),
    .S(_04185_),
    .X(_04191_));
 sky130_fd_sc_hd__clkbuf_1 _18295_ (.A(_04191_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _18296_ (.A0(_04025_),
    .A1(\cur_mb_mem[232][6] ),
    .S(_04185_),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _18297_ (.A(_04192_),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_1 _18298_ (.A0(_04027_),
    .A1(\cur_mb_mem[232][7] ),
    .S(_04185_),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_1 _18299_ (.A(_04193_),
    .X(_02014_));
 sky130_fd_sc_hd__and3_1 _18300_ (.A(_08978_),
    .B(_04107_),
    .C(_04135_),
    .X(_04194_));
 sky130_fd_sc_hd__clkbuf_4 _18301_ (.A(_04194_),
    .X(_04195_));
 sky130_fd_sc_hd__mux2_1 _18302_ (.A0(net1718),
    .A1(_04049_),
    .S(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_1 _18303_ (.A(_04196_),
    .X(_02015_));
 sky130_fd_sc_hd__mux2_1 _18304_ (.A0(net1737),
    .A1(_04053_),
    .S(_04195_),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_1 _18305_ (.A(_04197_),
    .X(_02016_));
 sky130_fd_sc_hd__mux2_1 _18306_ (.A0(net1836),
    .A1(_04055_),
    .S(_04195_),
    .X(_04198_));
 sky130_fd_sc_hd__clkbuf_1 _18307_ (.A(_04198_),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _18308_ (.A0(net1805),
    .A1(_04057_),
    .S(_04195_),
    .X(_04199_));
 sky130_fd_sc_hd__clkbuf_1 _18309_ (.A(_04199_),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _18310_ (.A0(net922),
    .A1(_04059_),
    .S(_04195_),
    .X(_04200_));
 sky130_fd_sc_hd__clkbuf_1 _18311_ (.A(_04200_),
    .X(_02019_));
 sky130_fd_sc_hd__mux2_1 _18312_ (.A0(net1631),
    .A1(_04061_),
    .S(_04195_),
    .X(_04201_));
 sky130_fd_sc_hd__clkbuf_1 _18313_ (.A(_04201_),
    .X(_02020_));
 sky130_fd_sc_hd__mux2_1 _18314_ (.A0(net836),
    .A1(_04063_),
    .S(_04195_),
    .X(_04202_));
 sky130_fd_sc_hd__clkbuf_1 _18315_ (.A(_04202_),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_1 _18316_ (.A0(\cur_mb_mem[233][7] ),
    .A1(_04065_),
    .S(_04195_),
    .X(_04203_));
 sky130_fd_sc_hd__clkbuf_1 _18317_ (.A(_04203_),
    .X(_02022_));
 sky130_fd_sc_hd__clkbuf_4 _18318_ (.A(_08530_),
    .X(_04204_));
 sky130_fd_sc_hd__and3_1 _18319_ (.A(_02353_),
    .B(_04107_),
    .C(_04135_),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_4 _18320_ (.A(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__mux2_1 _18321_ (.A0(net1881),
    .A1(_04204_),
    .S(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_1 _18322_ (.A(_04207_),
    .X(_02023_));
 sky130_fd_sc_hd__buf_4 _18323_ (.A(_08535_),
    .X(_04208_));
 sky130_fd_sc_hd__mux2_1 _18324_ (.A0(net1887),
    .A1(_04208_),
    .S(_04206_),
    .X(_04209_));
 sky130_fd_sc_hd__clkbuf_1 _18325_ (.A(_04209_),
    .X(_02024_));
 sky130_fd_sc_hd__buf_4 _18326_ (.A(_08538_),
    .X(_04210_));
 sky130_fd_sc_hd__mux2_1 _18327_ (.A0(\cur_mb_mem[234][2] ),
    .A1(_04210_),
    .S(_04206_),
    .X(_04211_));
 sky130_fd_sc_hd__clkbuf_1 _18328_ (.A(_04211_),
    .X(_02025_));
 sky130_fd_sc_hd__clkbuf_4 _18329_ (.A(_08541_),
    .X(_04212_));
 sky130_fd_sc_hd__mux2_1 _18330_ (.A0(net1798),
    .A1(_04212_),
    .S(_04206_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_1 _18331_ (.A(_04213_),
    .X(_02026_));
 sky130_fd_sc_hd__buf_4 _18332_ (.A(_08544_),
    .X(_04214_));
 sky130_fd_sc_hd__mux2_1 _18333_ (.A0(net1907),
    .A1(_04214_),
    .S(_04206_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_1 _18334_ (.A(_04215_),
    .X(_02027_));
 sky130_fd_sc_hd__buf_4 _18335_ (.A(_08547_),
    .X(_04216_));
 sky130_fd_sc_hd__mux2_1 _18336_ (.A0(net1846),
    .A1(_04216_),
    .S(_04206_),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _18337_ (.A(_04217_),
    .X(_02028_));
 sky130_fd_sc_hd__clkbuf_4 _18338_ (.A(_08550_),
    .X(_04218_));
 sky130_fd_sc_hd__mux2_1 _18339_ (.A0(net1871),
    .A1(_04218_),
    .S(_04206_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _18340_ (.A(_04219_),
    .X(_02029_));
 sky130_fd_sc_hd__buf_2 _18341_ (.A(_08553_),
    .X(_04220_));
 sky130_fd_sc_hd__mux2_1 _18342_ (.A0(\cur_mb_mem[234][7] ),
    .A1(_04220_),
    .S(_04206_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_1 _18343_ (.A(_04221_),
    .X(_02030_));
 sky130_fd_sc_hd__and3_1 _18344_ (.A(_02526_),
    .B(_04107_),
    .C(_04135_),
    .X(_04222_));
 sky130_fd_sc_hd__buf_4 _18345_ (.A(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__mux2_1 _18346_ (.A0(\cur_mb_mem[235][0] ),
    .A1(_04204_),
    .S(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_1 _18347_ (.A(_04224_),
    .X(_02031_));
 sky130_fd_sc_hd__mux2_1 _18348_ (.A0(\cur_mb_mem[235][1] ),
    .A1(_04208_),
    .S(_04223_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_1 _18349_ (.A(_04225_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _18350_ (.A0(\cur_mb_mem[235][2] ),
    .A1(_04210_),
    .S(_04223_),
    .X(_04226_));
 sky130_fd_sc_hd__clkbuf_1 _18351_ (.A(_04226_),
    .X(_02033_));
 sky130_fd_sc_hd__mux2_1 _18352_ (.A0(\cur_mb_mem[235][3] ),
    .A1(_04212_),
    .S(_04223_),
    .X(_04227_));
 sky130_fd_sc_hd__clkbuf_1 _18353_ (.A(_04227_),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _18354_ (.A0(net1908),
    .A1(_04214_),
    .S(_04223_),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_1 _18355_ (.A(_04228_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _18356_ (.A0(net1875),
    .A1(_04216_),
    .S(_04223_),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_1 _18357_ (.A(_04229_),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _18358_ (.A0(net1703),
    .A1(_04218_),
    .S(_04223_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_1 _18359_ (.A(_04230_),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _18360_ (.A0(net1716),
    .A1(_04220_),
    .S(_04223_),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _18361_ (.A(_04231_),
    .X(_02038_));
 sky130_fd_sc_hd__and3_1 _18362_ (.A(_02374_),
    .B(_04107_),
    .C(_04135_),
    .X(_04232_));
 sky130_fd_sc_hd__buf_4 _18363_ (.A(_04232_),
    .X(_04233_));
 sky130_fd_sc_hd__mux2_1 _18364_ (.A0(\cur_mb_mem[236][0] ),
    .A1(_04204_),
    .S(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__clkbuf_1 _18365_ (.A(_04234_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _18366_ (.A0(net1629),
    .A1(_04208_),
    .S(_04233_),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _18367_ (.A(_04235_),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _18368_ (.A0(net1857),
    .A1(_04210_),
    .S(_04233_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_1 _18369_ (.A(_04236_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _18370_ (.A0(net1876),
    .A1(_04212_),
    .S(_04233_),
    .X(_04237_));
 sky130_fd_sc_hd__clkbuf_1 _18371_ (.A(_04237_),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _18372_ (.A0(net1151),
    .A1(_04214_),
    .S(_04233_),
    .X(_04238_));
 sky130_fd_sc_hd__clkbuf_1 _18373_ (.A(_04238_),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_1 _18374_ (.A0(net640),
    .A1(_04216_),
    .S(_04233_),
    .X(_04239_));
 sky130_fd_sc_hd__clkbuf_1 _18375_ (.A(_04239_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _18376_ (.A0(net1824),
    .A1(_04218_),
    .S(_04233_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_1 _18377_ (.A(_04240_),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _18378_ (.A0(net1658),
    .A1(_04220_),
    .S(_04233_),
    .X(_04241_));
 sky130_fd_sc_hd__clkbuf_1 _18379_ (.A(_04241_),
    .X(_02046_));
 sky130_fd_sc_hd__and3_1 _18380_ (.A(_09025_),
    .B(_06067_),
    .C(_04135_),
    .X(_04242_));
 sky130_fd_sc_hd__buf_4 _18381_ (.A(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__mux2_1 _18382_ (.A0(net814),
    .A1(_04204_),
    .S(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _18383_ (.A(_04244_),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _18384_ (.A0(\cur_mb_mem[237][1] ),
    .A1(_04208_),
    .S(_04243_),
    .X(_04245_));
 sky130_fd_sc_hd__clkbuf_1 _18385_ (.A(_04245_),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _18386_ (.A0(net1822),
    .A1(_04210_),
    .S(_04243_),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_1 _18387_ (.A(_04246_),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _18388_ (.A0(net1931),
    .A1(_04212_),
    .S(_04243_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_1 _18389_ (.A(_04247_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _18390_ (.A0(net367),
    .A1(_04214_),
    .S(_04243_),
    .X(_04248_));
 sky130_fd_sc_hd__clkbuf_1 _18391_ (.A(_04248_),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _18392_ (.A0(net706),
    .A1(_04216_),
    .S(_04243_),
    .X(_04249_));
 sky130_fd_sc_hd__clkbuf_1 _18393_ (.A(_04249_),
    .X(_02052_));
 sky130_fd_sc_hd__mux2_1 _18394_ (.A0(net1912),
    .A1(_04218_),
    .S(_04243_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_1 _18395_ (.A(_04250_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _18396_ (.A0(\cur_mb_mem[237][7] ),
    .A1(_04220_),
    .S(_04243_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_1 _18397_ (.A(_04251_),
    .X(_02054_));
 sky130_fd_sc_hd__and3_1 _18398_ (.A(_09036_),
    .B(_06067_),
    .C(_04135_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_4 _18399_ (.A(_04252_),
    .X(_04253_));
 sky130_fd_sc_hd__mux2_1 _18400_ (.A0(net1893),
    .A1(_04204_),
    .S(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__clkbuf_1 _18401_ (.A(_04254_),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_1 _18402_ (.A0(net1677),
    .A1(_04208_),
    .S(_04253_),
    .X(_04255_));
 sky130_fd_sc_hd__clkbuf_1 _18403_ (.A(_04255_),
    .X(_02056_));
 sky130_fd_sc_hd__mux2_1 _18404_ (.A0(net1664),
    .A1(_04210_),
    .S(_04253_),
    .X(_04256_));
 sky130_fd_sc_hd__clkbuf_1 _18405_ (.A(_04256_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _18406_ (.A0(net1898),
    .A1(_04212_),
    .S(_04253_),
    .X(_04257_));
 sky130_fd_sc_hd__clkbuf_1 _18407_ (.A(_04257_),
    .X(_02058_));
 sky130_fd_sc_hd__mux2_1 _18408_ (.A0(net1145),
    .A1(_04214_),
    .S(_04253_),
    .X(_04258_));
 sky130_fd_sc_hd__clkbuf_1 _18409_ (.A(_04258_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _18410_ (.A0(net1525),
    .A1(_04216_),
    .S(_04253_),
    .X(_04259_));
 sky130_fd_sc_hd__clkbuf_1 _18411_ (.A(_04259_),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_1 _18412_ (.A0(net1785),
    .A1(_04218_),
    .S(_04253_),
    .X(_04260_));
 sky130_fd_sc_hd__clkbuf_1 _18413_ (.A(_04260_),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _18414_ (.A0(net1666),
    .A1(_04220_),
    .S(_04253_),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_1 _18415_ (.A(_04261_),
    .X(_02062_));
 sky130_fd_sc_hd__clkbuf_4 _18416_ (.A(_08880_),
    .X(_04262_));
 sky130_fd_sc_hd__and3_1 _18417_ (.A(_02406_),
    .B(_06067_),
    .C(_04262_),
    .X(_04263_));
 sky130_fd_sc_hd__buf_4 _18418_ (.A(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__mux2_1 _18419_ (.A0(\cur_mb_mem[239][0] ),
    .A1(_04204_),
    .S(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _18420_ (.A(_04265_),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_1 _18421_ (.A0(\cur_mb_mem[239][1] ),
    .A1(_04208_),
    .S(_04264_),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_1 _18422_ (.A(_04266_),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _18423_ (.A0(net1914),
    .A1(_04210_),
    .S(_04264_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_1 _18424_ (.A(_04267_),
    .X(_02065_));
 sky130_fd_sc_hd__mux2_1 _18425_ (.A0(\cur_mb_mem[239][3] ),
    .A1(_04212_),
    .S(_04264_),
    .X(_04268_));
 sky130_fd_sc_hd__clkbuf_1 _18426_ (.A(_04268_),
    .X(_02066_));
 sky130_fd_sc_hd__mux2_1 _18427_ (.A0(\cur_mb_mem[239][4] ),
    .A1(_04214_),
    .S(_04264_),
    .X(_04269_));
 sky130_fd_sc_hd__clkbuf_1 _18428_ (.A(_04269_),
    .X(_02067_));
 sky130_fd_sc_hd__mux2_1 _18429_ (.A0(\cur_mb_mem[239][5] ),
    .A1(_04216_),
    .S(_04264_),
    .X(_04270_));
 sky130_fd_sc_hd__clkbuf_1 _18430_ (.A(_04270_),
    .X(_02068_));
 sky130_fd_sc_hd__mux2_1 _18431_ (.A0(\cur_mb_mem[239][6] ),
    .A1(_04218_),
    .S(_04264_),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_1 _18432_ (.A(_04271_),
    .X(_02069_));
 sky130_fd_sc_hd__mux2_1 _18433_ (.A0(\cur_mb_mem[239][7] ),
    .A1(_04220_),
    .S(_04264_),
    .X(_04272_));
 sky130_fd_sc_hd__clkbuf_1 _18434_ (.A(_04272_),
    .X(_02070_));
 sky130_fd_sc_hd__buf_4 _18435_ (.A(_04432_),
    .X(_04273_));
 sky130_fd_sc_hd__nand2_8 _18436_ (.A(_04273_),
    .B(_08882_),
    .Y(_04274_));
 sky130_fd_sc_hd__mux2_1 _18437_ (.A0(_04012_),
    .A1(\cur_mb_mem[240][0] ),
    .S(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__clkbuf_1 _18438_ (.A(_04275_),
    .X(_02071_));
 sky130_fd_sc_hd__mux2_1 _18439_ (.A0(_04015_),
    .A1(net1840),
    .S(_04274_),
    .X(_04276_));
 sky130_fd_sc_hd__clkbuf_1 _18440_ (.A(_04276_),
    .X(_02072_));
 sky130_fd_sc_hd__mux2_1 _18441_ (.A0(_04017_),
    .A1(net702),
    .S(_04274_),
    .X(_04277_));
 sky130_fd_sc_hd__clkbuf_1 _18442_ (.A(_04277_),
    .X(_02073_));
 sky130_fd_sc_hd__mux2_1 _18443_ (.A0(_04019_),
    .A1(net1984),
    .S(_04274_),
    .X(_04278_));
 sky130_fd_sc_hd__clkbuf_1 _18444_ (.A(_04278_),
    .X(_02074_));
 sky130_fd_sc_hd__mux2_1 _18445_ (.A0(_04021_),
    .A1(net1812),
    .S(_04274_),
    .X(_04279_));
 sky130_fd_sc_hd__clkbuf_1 _18446_ (.A(_04279_),
    .X(_02075_));
 sky130_fd_sc_hd__mux2_1 _18447_ (.A0(_04023_),
    .A1(net1796),
    .S(_04274_),
    .X(_04280_));
 sky130_fd_sc_hd__clkbuf_1 _18448_ (.A(_04280_),
    .X(_02076_));
 sky130_fd_sc_hd__mux2_1 _18449_ (.A0(_04025_),
    .A1(\cur_mb_mem[240][6] ),
    .S(_04274_),
    .X(_04281_));
 sky130_fd_sc_hd__clkbuf_1 _18450_ (.A(_04281_),
    .X(_02077_));
 sky130_fd_sc_hd__mux2_1 _18451_ (.A0(_04027_),
    .A1(\cur_mb_mem[240][7] ),
    .S(_04274_),
    .X(_04282_));
 sky130_fd_sc_hd__clkbuf_1 _18452_ (.A(_04282_),
    .X(_02078_));
 sky130_fd_sc_hd__or4_1 _18453_ (.A(_05213_),
    .B(_05160_),
    .C(_05963_),
    .D(_08532_),
    .X(_04283_));
 sky130_fd_sc_hd__buf_4 _18454_ (.A(_04283_),
    .X(_04284_));
 sky130_fd_sc_hd__mux2_1 _18455_ (.A0(_04012_),
    .A1(\cur_mb_mem[241][0] ),
    .S(_04284_),
    .X(_04285_));
 sky130_fd_sc_hd__clkbuf_1 _18456_ (.A(_04285_),
    .X(_02079_));
 sky130_fd_sc_hd__mux2_1 _18457_ (.A0(_04015_),
    .A1(\cur_mb_mem[241][1] ),
    .S(_04284_),
    .X(_04286_));
 sky130_fd_sc_hd__clkbuf_1 _18458_ (.A(_04286_),
    .X(_02080_));
 sky130_fd_sc_hd__mux2_1 _18459_ (.A0(_04017_),
    .A1(\cur_mb_mem[241][2] ),
    .S(_04284_),
    .X(_04287_));
 sky130_fd_sc_hd__clkbuf_1 _18460_ (.A(_04287_),
    .X(_02081_));
 sky130_fd_sc_hd__mux2_1 _18461_ (.A0(_04019_),
    .A1(net1755),
    .S(_04284_),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_1 _18462_ (.A(_04288_),
    .X(_02082_));
 sky130_fd_sc_hd__mux2_1 _18463_ (.A0(_04021_),
    .A1(net1795),
    .S(_04284_),
    .X(_04289_));
 sky130_fd_sc_hd__clkbuf_1 _18464_ (.A(_04289_),
    .X(_02083_));
 sky130_fd_sc_hd__mux2_1 _18465_ (.A0(_04023_),
    .A1(net1844),
    .S(_04284_),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_1 _18466_ (.A(_04290_),
    .X(_02084_));
 sky130_fd_sc_hd__mux2_1 _18467_ (.A0(_04025_),
    .A1(\cur_mb_mem[241][6] ),
    .S(_04284_),
    .X(_04291_));
 sky130_fd_sc_hd__clkbuf_1 _18468_ (.A(_04291_),
    .X(_02085_));
 sky130_fd_sc_hd__mux2_1 _18469_ (.A0(_04027_),
    .A1(\cur_mb_mem[241][7] ),
    .S(_04284_),
    .X(_04292_));
 sky130_fd_sc_hd__clkbuf_1 _18470_ (.A(_04292_),
    .X(_02086_));
 sky130_fd_sc_hd__nand2_4 _18471_ (.A(_06335_),
    .B(_08979_),
    .Y(_04293_));
 sky130_fd_sc_hd__mux2_1 _18472_ (.A0(_04012_),
    .A1(net1688),
    .S(_04293_),
    .X(_04294_));
 sky130_fd_sc_hd__clkbuf_1 _18473_ (.A(_04294_),
    .X(_02087_));
 sky130_fd_sc_hd__mux2_1 _18474_ (.A0(_04015_),
    .A1(\cur_mb_mem[242][1] ),
    .S(_04293_),
    .X(_04295_));
 sky130_fd_sc_hd__clkbuf_1 _18475_ (.A(_04295_),
    .X(_02088_));
 sky130_fd_sc_hd__mux2_1 _18476_ (.A0(_04017_),
    .A1(net1541),
    .S(_04293_),
    .X(_04296_));
 sky130_fd_sc_hd__clkbuf_1 _18477_ (.A(_04296_),
    .X(_02089_));
 sky130_fd_sc_hd__mux2_1 _18478_ (.A0(_04019_),
    .A1(\cur_mb_mem[242][3] ),
    .S(_04293_),
    .X(_04297_));
 sky130_fd_sc_hd__clkbuf_1 _18479_ (.A(_04297_),
    .X(_02090_));
 sky130_fd_sc_hd__mux2_1 _18480_ (.A0(_04021_),
    .A1(net1809),
    .S(_04293_),
    .X(_04298_));
 sky130_fd_sc_hd__clkbuf_1 _18481_ (.A(_04298_),
    .X(_02091_));
 sky130_fd_sc_hd__mux2_1 _18482_ (.A0(_04023_),
    .A1(net1761),
    .S(_04293_),
    .X(_04299_));
 sky130_fd_sc_hd__clkbuf_1 _18483_ (.A(_04299_),
    .X(_02092_));
 sky130_fd_sc_hd__mux2_1 _18484_ (.A0(_04025_),
    .A1(\cur_mb_mem[242][6] ),
    .S(_04293_),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _18485_ (.A(_04300_),
    .X(_02093_));
 sky130_fd_sc_hd__mux2_1 _18486_ (.A0(_04027_),
    .A1(\cur_mb_mem[242][7] ),
    .S(_04293_),
    .X(_04301_));
 sky130_fd_sc_hd__clkbuf_1 _18487_ (.A(_04301_),
    .X(_02094_));
 sky130_fd_sc_hd__and3_1 _18488_ (.A(_04273_),
    .B(_06064_),
    .C(_04262_),
    .X(_04302_));
 sky130_fd_sc_hd__buf_4 _18489_ (.A(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__mux2_1 _18490_ (.A0(net1470),
    .A1(_04204_),
    .S(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__clkbuf_1 _18491_ (.A(_04304_),
    .X(_02095_));
 sky130_fd_sc_hd__mux2_1 _18492_ (.A0(net1894),
    .A1(_04208_),
    .S(_04303_),
    .X(_04305_));
 sky130_fd_sc_hd__clkbuf_1 _18493_ (.A(_04305_),
    .X(_02096_));
 sky130_fd_sc_hd__mux2_1 _18494_ (.A0(\cur_mb_mem[243][2] ),
    .A1(_04210_),
    .S(_04303_),
    .X(_04306_));
 sky130_fd_sc_hd__clkbuf_1 _18495_ (.A(_04306_),
    .X(_02097_));
 sky130_fd_sc_hd__mux2_1 _18496_ (.A0(\cur_mb_mem[243][3] ),
    .A1(_04212_),
    .S(_04303_),
    .X(_04307_));
 sky130_fd_sc_hd__clkbuf_1 _18497_ (.A(_04307_),
    .X(_02098_));
 sky130_fd_sc_hd__mux2_1 _18498_ (.A0(net948),
    .A1(_04214_),
    .S(_04303_),
    .X(_04308_));
 sky130_fd_sc_hd__clkbuf_1 _18499_ (.A(_04308_),
    .X(_02099_));
 sky130_fd_sc_hd__mux2_1 _18500_ (.A0(net1384),
    .A1(_04216_),
    .S(_04303_),
    .X(_04309_));
 sky130_fd_sc_hd__clkbuf_1 _18501_ (.A(_04309_),
    .X(_02100_));
 sky130_fd_sc_hd__mux2_1 _18502_ (.A0(\cur_mb_mem[243][6] ),
    .A1(_04218_),
    .S(_04303_),
    .X(_04310_));
 sky130_fd_sc_hd__clkbuf_1 _18503_ (.A(_04310_),
    .X(_02101_));
 sky130_fd_sc_hd__mux2_1 _18504_ (.A0(\cur_mb_mem[243][7] ),
    .A1(_04220_),
    .S(_04303_),
    .X(_04311_));
 sky130_fd_sc_hd__clkbuf_1 _18505_ (.A(_04311_),
    .X(_02102_));
 sky130_fd_sc_hd__nand2_8 _18506_ (.A(_06167_),
    .B(_08979_),
    .Y(_04312_));
 sky130_fd_sc_hd__mux2_1 _18507_ (.A0(_04012_),
    .A1(net1967),
    .S(_04312_),
    .X(_04313_));
 sky130_fd_sc_hd__clkbuf_1 _18508_ (.A(_04313_),
    .X(_02103_));
 sky130_fd_sc_hd__mux2_1 _18509_ (.A0(_04015_),
    .A1(\cur_mb_mem[244][1] ),
    .S(_04312_),
    .X(_04314_));
 sky130_fd_sc_hd__clkbuf_1 _18510_ (.A(_04314_),
    .X(_02104_));
 sky130_fd_sc_hd__mux2_1 _18511_ (.A0(_04017_),
    .A1(\cur_mb_mem[244][2] ),
    .S(_04312_),
    .X(_04315_));
 sky130_fd_sc_hd__clkbuf_1 _18512_ (.A(_04315_),
    .X(_02105_));
 sky130_fd_sc_hd__mux2_1 _18513_ (.A0(_04019_),
    .A1(net771),
    .S(_04312_),
    .X(_04316_));
 sky130_fd_sc_hd__clkbuf_1 _18514_ (.A(_04316_),
    .X(_02106_));
 sky130_fd_sc_hd__mux2_1 _18515_ (.A0(_04021_),
    .A1(\cur_mb_mem[244][4] ),
    .S(_04312_),
    .X(_04317_));
 sky130_fd_sc_hd__clkbuf_1 _18516_ (.A(_04317_),
    .X(_02107_));
 sky130_fd_sc_hd__mux2_1 _18517_ (.A0(_04023_),
    .A1(\cur_mb_mem[244][5] ),
    .S(_04312_),
    .X(_04318_));
 sky130_fd_sc_hd__clkbuf_1 _18518_ (.A(_04318_),
    .X(_02108_));
 sky130_fd_sc_hd__mux2_1 _18519_ (.A0(_04025_),
    .A1(\cur_mb_mem[244][6] ),
    .S(_04312_),
    .X(_04319_));
 sky130_fd_sc_hd__clkbuf_1 _18520_ (.A(_04319_),
    .X(_02109_));
 sky130_fd_sc_hd__mux2_1 _18521_ (.A0(_04027_),
    .A1(\cur_mb_mem[244][7] ),
    .S(_04312_),
    .X(_04320_));
 sky130_fd_sc_hd__clkbuf_1 _18522_ (.A(_04320_),
    .X(_02110_));
 sky130_fd_sc_hd__and3_1 _18523_ (.A(_04273_),
    .B(_06133_),
    .C(_04262_),
    .X(_04321_));
 sky130_fd_sc_hd__buf_4 _18524_ (.A(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__mux2_1 _18525_ (.A0(\cur_mb_mem[245][0] ),
    .A1(_04204_),
    .S(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__clkbuf_1 _18526_ (.A(_04323_),
    .X(_02111_));
 sky130_fd_sc_hd__mux2_1 _18527_ (.A0(\cur_mb_mem[245][1] ),
    .A1(_04208_),
    .S(_04322_),
    .X(_04324_));
 sky130_fd_sc_hd__clkbuf_1 _18528_ (.A(_04324_),
    .X(_02112_));
 sky130_fd_sc_hd__mux2_1 _18529_ (.A0(\cur_mb_mem[245][2] ),
    .A1(_04210_),
    .S(_04322_),
    .X(_04325_));
 sky130_fd_sc_hd__clkbuf_1 _18530_ (.A(_04325_),
    .X(_02113_));
 sky130_fd_sc_hd__mux2_1 _18531_ (.A0(net1989),
    .A1(_04212_),
    .S(_04322_),
    .X(_04326_));
 sky130_fd_sc_hd__clkbuf_1 _18532_ (.A(_04326_),
    .X(_02114_));
 sky130_fd_sc_hd__mux2_1 _18533_ (.A0(net1882),
    .A1(_04214_),
    .S(_04322_),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_1 _18534_ (.A(_04327_),
    .X(_02115_));
 sky130_fd_sc_hd__mux2_1 _18535_ (.A0(\cur_mb_mem[245][5] ),
    .A1(_04216_),
    .S(_04322_),
    .X(_04328_));
 sky130_fd_sc_hd__clkbuf_1 _18536_ (.A(_04328_),
    .X(_02116_));
 sky130_fd_sc_hd__mux2_1 _18537_ (.A0(net1661),
    .A1(_04218_),
    .S(_04322_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _18538_ (.A(_04329_),
    .X(_02117_));
 sky130_fd_sc_hd__mux2_1 _18539_ (.A0(net1656),
    .A1(_04220_),
    .S(_04322_),
    .X(_04330_));
 sky130_fd_sc_hd__clkbuf_1 _18540_ (.A(_04330_),
    .X(_02118_));
 sky130_fd_sc_hd__and3_1 _18541_ (.A(_04273_),
    .B(_06187_),
    .C(_04262_),
    .X(_04331_));
 sky130_fd_sc_hd__buf_4 _18542_ (.A(_04331_),
    .X(_04332_));
 sky130_fd_sc_hd__mux2_1 _18543_ (.A0(\cur_mb_mem[246][0] ),
    .A1(_04204_),
    .S(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__clkbuf_1 _18544_ (.A(_04333_),
    .X(_02119_));
 sky130_fd_sc_hd__mux2_1 _18545_ (.A0(\cur_mb_mem[246][1] ),
    .A1(_04208_),
    .S(_04332_),
    .X(_04334_));
 sky130_fd_sc_hd__clkbuf_1 _18546_ (.A(_04334_),
    .X(_02120_));
 sky130_fd_sc_hd__mux2_1 _18547_ (.A0(\cur_mb_mem[246][2] ),
    .A1(_04210_),
    .S(_04332_),
    .X(_04335_));
 sky130_fd_sc_hd__clkbuf_1 _18548_ (.A(_04335_),
    .X(_02121_));
 sky130_fd_sc_hd__mux2_1 _18549_ (.A0(net1762),
    .A1(_04212_),
    .S(_04332_),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_1 _18550_ (.A(_04336_),
    .X(_02122_));
 sky130_fd_sc_hd__mux2_1 _18551_ (.A0(\cur_mb_mem[246][4] ),
    .A1(_04214_),
    .S(_04332_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_1 _18552_ (.A(_04337_),
    .X(_02123_));
 sky130_fd_sc_hd__mux2_1 _18553_ (.A0(\cur_mb_mem[246][5] ),
    .A1(_04216_),
    .S(_04332_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_1 _18554_ (.A(_04338_),
    .X(_02124_));
 sky130_fd_sc_hd__mux2_1 _18555_ (.A0(\cur_mb_mem[246][6] ),
    .A1(_04218_),
    .S(_04332_),
    .X(_04339_));
 sky130_fd_sc_hd__clkbuf_1 _18556_ (.A(_04339_),
    .X(_02125_));
 sky130_fd_sc_hd__mux2_1 _18557_ (.A0(\cur_mb_mem[246][7] ),
    .A1(_04220_),
    .S(_04332_),
    .X(_04340_));
 sky130_fd_sc_hd__clkbuf_1 _18558_ (.A(_04340_),
    .X(_02126_));
 sky130_fd_sc_hd__and3_1 _18559_ (.A(_04273_),
    .B(_06103_),
    .C(_04262_),
    .X(_04341_));
 sky130_fd_sc_hd__buf_4 _18560_ (.A(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__mux2_1 _18561_ (.A0(net1700),
    .A1(_04204_),
    .S(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_1 _18562_ (.A(_04343_),
    .X(_02127_));
 sky130_fd_sc_hd__mux2_1 _18563_ (.A0(\cur_mb_mem[247][1] ),
    .A1(_04208_),
    .S(_04342_),
    .X(_04344_));
 sky130_fd_sc_hd__clkbuf_1 _18564_ (.A(_04344_),
    .X(_02128_));
 sky130_fd_sc_hd__mux2_1 _18565_ (.A0(net1817),
    .A1(_04210_),
    .S(_04342_),
    .X(_04345_));
 sky130_fd_sc_hd__clkbuf_1 _18566_ (.A(_04345_),
    .X(_02129_));
 sky130_fd_sc_hd__mux2_1 _18567_ (.A0(net1756),
    .A1(_04212_),
    .S(_04342_),
    .X(_04346_));
 sky130_fd_sc_hd__clkbuf_1 _18568_ (.A(_04346_),
    .X(_02130_));
 sky130_fd_sc_hd__mux2_1 _18569_ (.A0(net652),
    .A1(_04214_),
    .S(_04342_),
    .X(_04347_));
 sky130_fd_sc_hd__clkbuf_1 _18570_ (.A(_04347_),
    .X(_02131_));
 sky130_fd_sc_hd__mux2_1 _18571_ (.A0(net826),
    .A1(_04216_),
    .S(_04342_),
    .X(_04348_));
 sky130_fd_sc_hd__clkbuf_1 _18572_ (.A(_04348_),
    .X(_02132_));
 sky130_fd_sc_hd__mux2_1 _18573_ (.A0(\cur_mb_mem[247][6] ),
    .A1(_04218_),
    .S(_04342_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _18574_ (.A(_04349_),
    .X(_02133_));
 sky130_fd_sc_hd__mux2_1 _18575_ (.A0(net1905),
    .A1(_04220_),
    .S(_04342_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_1 _18576_ (.A(_04350_),
    .X(_02134_));
 sky130_fd_sc_hd__nand2_8 _18577_ (.A(_06411_),
    .B(_08979_),
    .Y(_04351_));
 sky130_fd_sc_hd__mux2_1 _18578_ (.A0(_08531_),
    .A1(net1381),
    .S(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_1 _18579_ (.A(_04352_),
    .X(_02135_));
 sky130_fd_sc_hd__mux2_1 _18580_ (.A0(_08536_),
    .A1(\cur_mb_mem[248][1] ),
    .S(_04351_),
    .X(_04353_));
 sky130_fd_sc_hd__clkbuf_1 _18581_ (.A(_04353_),
    .X(_02136_));
 sky130_fd_sc_hd__mux2_1 _18582_ (.A0(_08539_),
    .A1(net1544),
    .S(_04351_),
    .X(_04354_));
 sky130_fd_sc_hd__clkbuf_1 _18583_ (.A(_04354_),
    .X(_02137_));
 sky130_fd_sc_hd__mux2_1 _18584_ (.A0(_08542_),
    .A1(net1974),
    .S(_04351_),
    .X(_04355_));
 sky130_fd_sc_hd__clkbuf_1 _18585_ (.A(_04355_),
    .X(_02138_));
 sky130_fd_sc_hd__mux2_1 _18586_ (.A0(_08545_),
    .A1(net1458),
    .S(_04351_),
    .X(_04356_));
 sky130_fd_sc_hd__clkbuf_1 _18587_ (.A(_04356_),
    .X(_02139_));
 sky130_fd_sc_hd__mux2_1 _18588_ (.A0(_08548_),
    .A1(net1417),
    .S(_04351_),
    .X(_04357_));
 sky130_fd_sc_hd__clkbuf_1 _18589_ (.A(_04357_),
    .X(_02140_));
 sky130_fd_sc_hd__mux2_1 _18590_ (.A0(_08551_),
    .A1(net1374),
    .S(_04351_),
    .X(_04358_));
 sky130_fd_sc_hd__clkbuf_1 _18591_ (.A(_04358_),
    .X(_02141_));
 sky130_fd_sc_hd__mux2_1 _18592_ (.A0(_08554_),
    .A1(net1149),
    .S(_04351_),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_1 _18593_ (.A(_04359_),
    .X(_02142_));
 sky130_fd_sc_hd__and3_1 _18594_ (.A(_04273_),
    .B(_05912_),
    .C(_04262_),
    .X(_04360_));
 sky130_fd_sc_hd__buf_6 _18595_ (.A(_04360_),
    .X(_04361_));
 sky130_fd_sc_hd__mux2_1 _18596_ (.A0(net433),
    .A1(_02327_),
    .S(_04361_),
    .X(_04362_));
 sky130_fd_sc_hd__clkbuf_1 _18597_ (.A(_04362_),
    .X(_02143_));
 sky130_fd_sc_hd__mux2_1 _18598_ (.A0(\cur_mb_mem[249][1] ),
    .A1(_02332_),
    .S(_04361_),
    .X(_04363_));
 sky130_fd_sc_hd__clkbuf_1 _18599_ (.A(_04363_),
    .X(_02144_));
 sky130_fd_sc_hd__mux2_1 _18600_ (.A0(net598),
    .A1(_02335_),
    .S(_04361_),
    .X(_04364_));
 sky130_fd_sc_hd__clkbuf_1 _18601_ (.A(_04364_),
    .X(_02145_));
 sky130_fd_sc_hd__mux2_1 _18602_ (.A0(net405),
    .A1(_02338_),
    .S(_04361_),
    .X(_04365_));
 sky130_fd_sc_hd__clkbuf_1 _18603_ (.A(_04365_),
    .X(_02146_));
 sky130_fd_sc_hd__mux2_1 _18604_ (.A0(net957),
    .A1(_02341_),
    .S(_04361_),
    .X(_04366_));
 sky130_fd_sc_hd__clkbuf_1 _18605_ (.A(_04366_),
    .X(_02147_));
 sky130_fd_sc_hd__mux2_1 _18606_ (.A0(net583),
    .A1(_02344_),
    .S(_04361_),
    .X(_04367_));
 sky130_fd_sc_hd__clkbuf_1 _18607_ (.A(_04367_),
    .X(_02148_));
 sky130_fd_sc_hd__mux2_1 _18608_ (.A0(net1654),
    .A1(_02347_),
    .S(_04361_),
    .X(_04368_));
 sky130_fd_sc_hd__clkbuf_1 _18609_ (.A(_04368_),
    .X(_02149_));
 sky130_fd_sc_hd__mux2_1 _18610_ (.A0(net1316),
    .A1(_02350_),
    .S(_04361_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_1 _18611_ (.A(_04369_),
    .X(_02150_));
 sky130_fd_sc_hd__and3_1 _18612_ (.A(_04273_),
    .B(_06035_),
    .C(_04262_),
    .X(_04370_));
 sky130_fd_sc_hd__clkbuf_8 _18613_ (.A(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__mux2_1 _18614_ (.A0(net1035),
    .A1(_02327_),
    .S(_04371_),
    .X(_04372_));
 sky130_fd_sc_hd__clkbuf_1 _18615_ (.A(_04372_),
    .X(_02151_));
 sky130_fd_sc_hd__mux2_1 _18616_ (.A0(net1478),
    .A1(_02332_),
    .S(_04371_),
    .X(_04373_));
 sky130_fd_sc_hd__clkbuf_1 _18617_ (.A(_04373_),
    .X(_02152_));
 sky130_fd_sc_hd__mux2_1 _18618_ (.A0(net1270),
    .A1(_02335_),
    .S(_04371_),
    .X(_04374_));
 sky130_fd_sc_hd__clkbuf_1 _18619_ (.A(_04374_),
    .X(_02153_));
 sky130_fd_sc_hd__mux2_1 _18620_ (.A0(net1422),
    .A1(_02338_),
    .S(_04371_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_1 _18621_ (.A(_04375_),
    .X(_02154_));
 sky130_fd_sc_hd__mux2_1 _18622_ (.A0(net1528),
    .A1(_02341_),
    .S(_04371_),
    .X(_04376_));
 sky130_fd_sc_hd__clkbuf_1 _18623_ (.A(_04376_),
    .X(_02155_));
 sky130_fd_sc_hd__mux2_1 _18624_ (.A0(net797),
    .A1(_02344_),
    .S(_04371_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_1 _18625_ (.A(_04377_),
    .X(_02156_));
 sky130_fd_sc_hd__mux2_1 _18626_ (.A0(net1830),
    .A1(_02347_),
    .S(_04371_),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_1 _18627_ (.A(_04378_),
    .X(_02157_));
 sky130_fd_sc_hd__mux2_1 _18628_ (.A0(net1074),
    .A1(_02350_),
    .S(_04371_),
    .X(_04379_));
 sky130_fd_sc_hd__clkbuf_1 _18629_ (.A(_04379_),
    .X(_02158_));
 sky130_fd_sc_hd__and3_1 _18630_ (.A(_04273_),
    .B(_06049_),
    .C(_04262_),
    .X(_04380_));
 sky130_fd_sc_hd__clkbuf_8 _18631_ (.A(_04380_),
    .X(_04381_));
 sky130_fd_sc_hd__mux2_1 _18632_ (.A0(net538),
    .A1(_02327_),
    .S(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__clkbuf_1 _18633_ (.A(_04382_),
    .X(_02159_));
 sky130_fd_sc_hd__mux2_1 _18634_ (.A0(net1326),
    .A1(_02332_),
    .S(_04381_),
    .X(_04383_));
 sky130_fd_sc_hd__clkbuf_1 _18635_ (.A(_04383_),
    .X(_02160_));
 sky130_fd_sc_hd__mux2_1 _18636_ (.A0(net729),
    .A1(_02335_),
    .S(_04381_),
    .X(_04384_));
 sky130_fd_sc_hd__clkbuf_1 _18637_ (.A(_04384_),
    .X(_02161_));
 sky130_fd_sc_hd__mux2_1 _18638_ (.A0(net611),
    .A1(_02338_),
    .S(_04381_),
    .X(_04385_));
 sky130_fd_sc_hd__clkbuf_1 _18639_ (.A(_04385_),
    .X(_02162_));
 sky130_fd_sc_hd__mux2_1 _18640_ (.A0(net420),
    .A1(_02341_),
    .S(_04381_),
    .X(_04386_));
 sky130_fd_sc_hd__clkbuf_1 _18641_ (.A(_04386_),
    .X(_02163_));
 sky130_fd_sc_hd__mux2_1 _18642_ (.A0(net1046),
    .A1(_02344_),
    .S(_04381_),
    .X(_04387_));
 sky130_fd_sc_hd__clkbuf_1 _18643_ (.A(_04387_),
    .X(_02164_));
 sky130_fd_sc_hd__mux2_1 _18644_ (.A0(net1577),
    .A1(_02347_),
    .S(_04381_),
    .X(_04388_));
 sky130_fd_sc_hd__clkbuf_1 _18645_ (.A(_04388_),
    .X(_02165_));
 sky130_fd_sc_hd__mux2_1 _18646_ (.A0(net1104),
    .A1(_02350_),
    .S(_04381_),
    .X(_04389_));
 sky130_fd_sc_hd__clkbuf_1 _18647_ (.A(_04389_),
    .X(_02166_));
 sky130_fd_sc_hd__and3_1 _18648_ (.A(_04273_),
    .B(_05989_),
    .C(_04262_),
    .X(_04390_));
 sky130_fd_sc_hd__clkbuf_8 _18649_ (.A(_04390_),
    .X(_04391_));
 sky130_fd_sc_hd__mux2_1 _18650_ (.A0(net609),
    .A1(_02327_),
    .S(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__clkbuf_1 _18651_ (.A(_04392_),
    .X(_02167_));
 sky130_fd_sc_hd__mux2_1 _18652_ (.A0(net384),
    .A1(_02332_),
    .S(_04391_),
    .X(_04393_));
 sky130_fd_sc_hd__clkbuf_1 _18653_ (.A(_04393_),
    .X(_02168_));
 sky130_fd_sc_hd__mux2_1 _18654_ (.A0(net338),
    .A1(_02335_),
    .S(_04391_),
    .X(_04394_));
 sky130_fd_sc_hd__clkbuf_1 _18655_ (.A(_04394_),
    .X(_02169_));
 sky130_fd_sc_hd__mux2_1 _18656_ (.A0(net1068),
    .A1(_02338_),
    .S(_04391_),
    .X(_04395_));
 sky130_fd_sc_hd__clkbuf_1 _18657_ (.A(_04395_),
    .X(_02170_));
 sky130_fd_sc_hd__mux2_1 _18658_ (.A0(net470),
    .A1(_02341_),
    .S(_04391_),
    .X(_04396_));
 sky130_fd_sc_hd__clkbuf_1 _18659_ (.A(_04396_),
    .X(_02171_));
 sky130_fd_sc_hd__mux2_1 _18660_ (.A0(net337),
    .A1(_02344_),
    .S(_04391_),
    .X(_04397_));
 sky130_fd_sc_hd__clkbuf_1 _18661_ (.A(_04397_),
    .X(_02172_));
 sky130_fd_sc_hd__mux2_1 _18662_ (.A0(net1307),
    .A1(_02347_),
    .S(_04391_),
    .X(_04398_));
 sky130_fd_sc_hd__clkbuf_1 _18663_ (.A(_04398_),
    .X(_02173_));
 sky130_fd_sc_hd__mux2_1 _18664_ (.A0(net1639),
    .A1(_02350_),
    .S(_04391_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_1 _18665_ (.A(_04399_),
    .X(_02174_));
 sky130_fd_sc_hd__and3_1 _18666_ (.A(_04273_),
    .B(_05961_),
    .C(_04262_),
    .X(_04400_));
 sky130_fd_sc_hd__buf_4 _18667_ (.A(_04400_),
    .X(_04401_));
 sky130_fd_sc_hd__mux2_1 _18668_ (.A0(net1633),
    .A1(_02327_),
    .S(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_1 _18669_ (.A(_04402_),
    .X(_02175_));
 sky130_fd_sc_hd__mux2_1 _18670_ (.A0(net1162),
    .A1(_02332_),
    .S(_04401_),
    .X(_04403_));
 sky130_fd_sc_hd__clkbuf_1 _18671_ (.A(_04403_),
    .X(_02176_));
 sky130_fd_sc_hd__mux2_1 _18672_ (.A0(net1750),
    .A1(_02335_),
    .S(_04401_),
    .X(_04404_));
 sky130_fd_sc_hd__clkbuf_1 _18673_ (.A(_04404_),
    .X(_02177_));
 sky130_fd_sc_hd__mux2_1 _18674_ (.A0(net1690),
    .A1(_02338_),
    .S(_04401_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_1 _18675_ (.A(_04405_),
    .X(_02178_));
 sky130_fd_sc_hd__mux2_1 _18676_ (.A0(net946),
    .A1(_02341_),
    .S(_04401_),
    .X(_04406_));
 sky130_fd_sc_hd__clkbuf_1 _18677_ (.A(_04406_),
    .X(_02179_));
 sky130_fd_sc_hd__mux2_1 _18678_ (.A0(net1223),
    .A1(_02344_),
    .S(_04401_),
    .X(_04407_));
 sky130_fd_sc_hd__clkbuf_1 _18679_ (.A(_04407_),
    .X(_02180_));
 sky130_fd_sc_hd__mux2_1 _18680_ (.A0(net894),
    .A1(_02347_),
    .S(_04401_),
    .X(_04408_));
 sky130_fd_sc_hd__clkbuf_1 _18681_ (.A(_04408_),
    .X(_02181_));
 sky130_fd_sc_hd__mux2_1 _18682_ (.A0(net959),
    .A1(_02350_),
    .S(_04401_),
    .X(_04409_));
 sky130_fd_sc_hd__clkbuf_1 _18683_ (.A(_04409_),
    .X(_02182_));
 sky130_fd_sc_hd__and3_1 _18684_ (.A(_04432_),
    .B(_06025_),
    .C(_08900_),
    .X(_04410_));
 sky130_fd_sc_hd__buf_6 _18685_ (.A(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__mux2_1 _18686_ (.A0(net589),
    .A1(_02327_),
    .S(_04411_),
    .X(_04412_));
 sky130_fd_sc_hd__clkbuf_1 _18687_ (.A(_04412_),
    .X(_02183_));
 sky130_fd_sc_hd__mux2_1 _18688_ (.A0(\cur_mb_mem[254][1] ),
    .A1(_02332_),
    .S(_04411_),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_1 _18689_ (.A(_04413_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _18690_ (.A0(net365),
    .A1(_02335_),
    .S(_04411_),
    .X(_04414_));
 sky130_fd_sc_hd__clkbuf_1 _18691_ (.A(_04414_),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_1 _18692_ (.A0(net432),
    .A1(_02338_),
    .S(_04411_),
    .X(_04415_));
 sky130_fd_sc_hd__clkbuf_1 _18693_ (.A(_04415_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _18694_ (.A0(net777),
    .A1(_02341_),
    .S(_04411_),
    .X(_04416_));
 sky130_fd_sc_hd__clkbuf_1 _18695_ (.A(_04416_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_1 _18696_ (.A0(net1089),
    .A1(_02344_),
    .S(_04411_),
    .X(_04417_));
 sky130_fd_sc_hd__clkbuf_1 _18697_ (.A(_04417_),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_1 _18698_ (.A0(net756),
    .A1(_02347_),
    .S(_04411_),
    .X(_04418_));
 sky130_fd_sc_hd__clkbuf_1 _18699_ (.A(_04418_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _18700_ (.A0(net1181),
    .A1(_02350_),
    .S(_04411_),
    .X(_04419_));
 sky130_fd_sc_hd__clkbuf_1 _18701_ (.A(_04419_),
    .X(_02190_));
 sky130_fd_sc_hd__dfxtp_1 _18702_ (.CLK(clknet_leaf_202_clk),
    .D(_00008_),
    .Q(\best_cand_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18703_ (.CLK(clknet_leaf_203_clk),
    .D(_00009_),
    .Q(\best_cand_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18704_ (.CLK(clknet_leaf_202_clk),
    .D(_00010_),
    .Q(\best_cand_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18705_ (.CLK(clknet_leaf_218_clk),
    .D(_00011_),
    .Q(\best_cand_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18706_ (.CLK(clknet_leaf_215_clk),
    .D(_00012_),
    .Q(\best_cand_x[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18707_ (.CLK(clknet_leaf_215_clk),
    .D(_00013_),
    .Q(\best_cand_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18708_ (.CLK(clknet_leaf_205_clk),
    .D(_00014_),
    .Q(\best_cand_x[6] ));
 sky130_fd_sc_hd__dfstp_1 _18709_ (.CLK(clknet_leaf_197_clk),
    .D(_00000_),
    .SET_B(net266),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _18710_ (.CLK(clknet_leaf_218_clk),
    .D(_00001_),
    .RESET_B(net266),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _18711_ (.CLK(clknet_leaf_217_clk),
    .D(_00003_),
    .RESET_B(net272),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _18712_ (.CLK(clknet_leaf_198_clk),
    .D(_00004_),
    .RESET_B(net266),
    .Q(\state[3] ));
 sky130_fd_sc_hd__dfrtp_4 _18713_ (.CLK(clknet_leaf_197_clk),
    .D(_00005_),
    .RESET_B(net266),
    .Q(\state[4] ));
 sky130_fd_sc_hd__dfrtp_2 _18714_ (.CLK(clknet_leaf_217_clk),
    .D(_00002_),
    .RESET_B(net272),
    .Q(\state[5] ));
 sky130_fd_sc_hd__dfrtp_4 _18715_ (.CLK(clknet_leaf_217_clk),
    .D(_00006_),
    .RESET_B(net272),
    .Q(\state[6] ));
 sky130_fd_sc_hd__dfrtp_2 _18716_ (.CLK(clknet_leaf_198_clk),
    .D(_00007_),
    .RESET_B(net266),
    .Q(\state[7] ));
 sky130_fd_sc_hd__dfstp_1 _18717_ (.CLK(clknet_leaf_189_clk),
    .D(_00015_),
    .SET_B(net268),
    .Q(\min_sad_reg[0] ));
 sky130_fd_sc_hd__dfstp_1 _18718_ (.CLK(clknet_leaf_188_clk),
    .D(_00016_),
    .SET_B(net268),
    .Q(\min_sad_reg[1] ));
 sky130_fd_sc_hd__dfstp_1 _18719_ (.CLK(clknet_leaf_189_clk),
    .D(_00017_),
    .SET_B(net269),
    .Q(\min_sad_reg[2] ));
 sky130_fd_sc_hd__dfstp_1 _18720_ (.CLK(clknet_leaf_188_clk),
    .D(_00018_),
    .SET_B(net269),
    .Q(\min_sad_reg[3] ));
 sky130_fd_sc_hd__dfstp_1 _18721_ (.CLK(clknet_leaf_188_clk),
    .D(_00019_),
    .SET_B(net269),
    .Q(\min_sad_reg[4] ));
 sky130_fd_sc_hd__dfstp_1 _18722_ (.CLK(clknet_leaf_187_clk),
    .D(_00020_),
    .SET_B(net269),
    .Q(\min_sad_reg[5] ));
 sky130_fd_sc_hd__dfstp_1 _18723_ (.CLK(clknet_leaf_187_clk),
    .D(_00021_),
    .SET_B(net269),
    .Q(\min_sad_reg[6] ));
 sky130_fd_sc_hd__dfstp_4 _18724_ (.CLK(clknet_leaf_190_clk),
    .D(_00022_),
    .SET_B(net268),
    .Q(\min_sad_reg[7] ));
 sky130_fd_sc_hd__dfstp_1 _18725_ (.CLK(clknet_leaf_190_clk),
    .D(_00023_),
    .SET_B(net268),
    .Q(\min_sad_reg[8] ));
 sky130_fd_sc_hd__dfstp_1 _18726_ (.CLK(clknet_leaf_190_clk),
    .D(_00024_),
    .SET_B(net268),
    .Q(\min_sad_reg[9] ));
 sky130_fd_sc_hd__dfstp_4 _18727_ (.CLK(clknet_leaf_200_clk),
    .D(_00025_),
    .SET_B(net270),
    .Q(\min_sad_reg[10] ));
 sky130_fd_sc_hd__dfstp_1 _18728_ (.CLK(clknet_leaf_190_clk),
    .D(_00026_),
    .SET_B(net268),
    .Q(\min_sad_reg[11] ));
 sky130_fd_sc_hd__dfstp_4 _18729_ (.CLK(clknet_leaf_190_clk),
    .D(_00027_),
    .SET_B(net268),
    .Q(\min_sad_reg[12] ));
 sky130_fd_sc_hd__dfstp_4 _18730_ (.CLK(clknet_leaf_194_clk),
    .D(_00028_),
    .SET_B(net267),
    .Q(\min_sad_reg[13] ));
 sky130_fd_sc_hd__dfstp_4 _18731_ (.CLK(clknet_leaf_194_clk),
    .D(_00029_),
    .SET_B(net267),
    .Q(\min_sad_reg[14] ));
 sky130_fd_sc_hd__dfstp_1 _18732_ (.CLK(clknet_leaf_197_clk),
    .D(_00030_),
    .SET_B(net266),
    .Q(\min_sad_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _18733_ (.CLK(clknet_leaf_256_clk),
    .D(_00031_),
    .Q(\cur_mb_mem[255][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18734_ (.CLK(clknet_leaf_273_clk),
    .D(_00032_),
    .Q(\cur_mb_mem[255][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18735_ (.CLK(clknet_leaf_255_clk),
    .D(_00033_),
    .Q(\cur_mb_mem[255][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18736_ (.CLK(clknet_leaf_257_clk),
    .D(_00034_),
    .Q(\cur_mb_mem[255][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18737_ (.CLK(clknet_leaf_273_clk),
    .D(_00035_),
    .Q(\cur_mb_mem[255][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18738_ (.CLK(clknet_leaf_273_clk),
    .D(_00036_),
    .Q(\cur_mb_mem[255][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18739_ (.CLK(clknet_leaf_318_clk),
    .D(_00037_),
    .Q(\cur_mb_mem[255][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18740_ (.CLK(clknet_leaf_237_clk),
    .D(_00038_),
    .Q(\cur_mb_mem[255][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18741_ (.CLK(clknet_leaf_199_clk),
    .D(_00039_),
    .Q(\best_point_idx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18742_ (.CLK(clknet_leaf_199_clk),
    .D(_00040_),
    .Q(\best_point_idx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18743_ (.CLK(clknet_leaf_199_clk),
    .D(_00041_),
    .Q(\best_point_idx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18744_ (.CLK(clknet_leaf_199_clk),
    .D(_00042_),
    .Q(\best_point_idx[3] ));
 sky130_fd_sc_hd__dfrtp_2 _18745_ (.CLK(clknet_leaf_206_clk),
    .D(_00043_),
    .RESET_B(net276),
    .Q(net172));
 sky130_fd_sc_hd__dfrtp_4 _18746_ (.CLK(clknet_leaf_200_clk),
    .D(_00044_),
    .RESET_B(net270),
    .Q(net173));
 sky130_fd_sc_hd__dfrtp_2 _18747_ (.CLK(clknet_leaf_201_clk),
    .D(_00045_),
    .RESET_B(net270),
    .Q(net174));
 sky130_fd_sc_hd__dfrtp_4 _18748_ (.CLK(clknet_leaf_218_clk),
    .D(_00046_),
    .RESET_B(net272),
    .Q(net175));
 sky130_fd_sc_hd__dfrtp_4 _18749_ (.CLK(clknet_leaf_215_clk),
    .D(_00047_),
    .RESET_B(net272),
    .Q(net176));
 sky130_fd_sc_hd__dfrtp_4 _18750_ (.CLK(clknet_5_30__leaf_clk),
    .D(_00048_),
    .RESET_B(net272),
    .Q(net177));
 sky130_fd_sc_hd__dfrtp_4 _18751_ (.CLK(clknet_leaf_202_clk),
    .D(_00049_),
    .RESET_B(net276),
    .Q(net178));
 sky130_fd_sc_hd__dfrtp_4 _18752_ (.CLK(clknet_leaf_212_clk),
    .D(_00050_),
    .RESET_B(net274),
    .Q(net179));
 sky130_fd_sc_hd__dfrtp_4 _18753_ (.CLK(clknet_leaf_206_clk),
    .D(_00051_),
    .RESET_B(net276),
    .Q(net180));
 sky130_fd_sc_hd__dfrtp_4 _18754_ (.CLK(clknet_leaf_196_clk),
    .D(_00052_),
    .RESET_B(net266),
    .Q(net181));
 sky130_fd_sc_hd__dfrtp_1 _18755_ (.CLK(clknet_leaf_211_clk),
    .D(_00053_),
    .RESET_B(net274),
    .Q(net182));
 sky130_fd_sc_hd__dfrtp_4 _18756_ (.CLK(clknet_leaf_196_clk),
    .D(_00054_),
    .RESET_B(net266),
    .Q(net183));
 sky130_fd_sc_hd__dfrtp_1 _18757_ (.CLK(clknet_leaf_202_clk),
    .D(_00055_),
    .RESET_B(net276),
    .Q(net184));
 sky130_fd_sc_hd__dfrtp_4 _18758_ (.CLK(clknet_leaf_202_clk),
    .D(_00056_),
    .RESET_B(net276),
    .Q(net191));
 sky130_fd_sc_hd__dfrtp_4 _18759_ (.CLK(clknet_leaf_190_clk),
    .D(_00057_),
    .RESET_B(net268),
    .Q(net192));
 sky130_fd_sc_hd__dfrtp_1 _18760_ (.CLK(clknet_leaf_188_clk),
    .D(_00058_),
    .RESET_B(net269),
    .Q(net193));
 sky130_fd_sc_hd__dfrtp_1 _18761_ (.CLK(clknet_leaf_188_clk),
    .D(_00059_),
    .RESET_B(net269),
    .Q(net194));
 sky130_fd_sc_hd__dfrtp_4 _18762_ (.CLK(clknet_leaf_187_clk),
    .D(_00060_),
    .RESET_B(net269),
    .Q(net195));
 sky130_fd_sc_hd__dfrtp_4 _18763_ (.CLK(clknet_leaf_187_clk),
    .D(_00061_),
    .RESET_B(net269),
    .Q(net196));
 sky130_fd_sc_hd__dfrtp_1 _18764_ (.CLK(clknet_leaf_291_clk),
    .D(_00062_),
    .RESET_B(net280),
    .Q(net197));
 sky130_fd_sc_hd__dfrtp_4 _18765_ (.CLK(clknet_leaf_191_clk),
    .D(_00063_),
    .RESET_B(net268),
    .Q(net198));
 sky130_fd_sc_hd__dfrtp_4 _18766_ (.CLK(clknet_leaf_191_clk),
    .D(_00064_),
    .RESET_B(net268),
    .Q(net199));
 sky130_fd_sc_hd__dfrtp_2 _18767_ (.CLK(clknet_leaf_276_clk),
    .D(_00065_),
    .RESET_B(net280),
    .Q(net185));
 sky130_fd_sc_hd__dfrtp_4 _18768_ (.CLK(clknet_leaf_193_clk),
    .D(_00066_),
    .RESET_B(net267),
    .Q(net186));
 sky130_fd_sc_hd__dfrtp_4 _18769_ (.CLK(clknet_leaf_284_clk),
    .D(_00067_),
    .RESET_B(net280),
    .Q(net187));
 sky130_fd_sc_hd__dfrtp_4 _18770_ (.CLK(clknet_leaf_291_clk),
    .D(_00068_),
    .RESET_B(net280),
    .Q(net188));
 sky130_fd_sc_hd__dfrtp_4 _18771_ (.CLK(clknet_leaf_291_clk),
    .D(_00069_),
    .RESET_B(net280),
    .Q(net189));
 sky130_fd_sc_hd__dfrtp_4 _18772_ (.CLK(clknet_leaf_197_clk),
    .D(_00070_),
    .RESET_B(net267),
    .Q(net190));
 sky130_fd_sc_hd__dfrtp_4 _18773_ (.CLK(clknet_leaf_201_clk),
    .D(_00071_),
    .RESET_B(net270),
    .Q(net139));
 sky130_fd_sc_hd__dfrtp_1 _18774_ (.CLK(clknet_leaf_202_clk),
    .D(_00072_),
    .RESET_B(net271),
    .Q(\center_x[0] ));
 sky130_fd_sc_hd__dfrtp_1 _18775_ (.CLK(clknet_leaf_201_clk),
    .D(_00073_),
    .RESET_B(net271),
    .Q(\center_x[1] ));
 sky130_fd_sc_hd__dfrtp_2 _18776_ (.CLK(clknet_leaf_202_clk),
    .D(_00074_),
    .RESET_B(net276),
    .Q(\center_x[2] ));
 sky130_fd_sc_hd__dfrtp_2 _18777_ (.CLK(clknet_leaf_217_clk),
    .D(_00075_),
    .RESET_B(net272),
    .Q(\center_x[3] ));
 sky130_fd_sc_hd__dfrtp_2 _18778_ (.CLK(clknet_leaf_215_clk),
    .D(_00076_),
    .RESET_B(net272),
    .Q(\center_x[4] ));
 sky130_fd_sc_hd__dfrtp_4 _18779_ (.CLK(clknet_leaf_215_clk),
    .D(_00077_),
    .RESET_B(net272),
    .Q(\center_x[5] ));
 sky130_fd_sc_hd__dfrtp_2 _18780_ (.CLK(clknet_leaf_206_clk),
    .D(_00078_),
    .RESET_B(net278),
    .Q(\center_x[6] ));
 sky130_fd_sc_hd__dfrtp_2 _18781_ (.CLK(clknet_leaf_202_clk),
    .D(_00079_),
    .RESET_B(net276),
    .Q(\center_y[0] ));
 sky130_fd_sc_hd__dfrtp_1 _18782_ (.CLK(clknet_leaf_217_clk),
    .D(net1570),
    .RESET_B(net273),
    .Q(\center_y[1] ));
 sky130_fd_sc_hd__dfrtp_4 _18783_ (.CLK(clknet_leaf_216_clk),
    .D(_00081_),
    .RESET_B(net274),
    .Q(\center_y[2] ));
 sky130_fd_sc_hd__dfrtp_2 _18784_ (.CLK(clknet_leaf_214_clk),
    .D(_00082_),
    .RESET_B(net274),
    .Q(\center_y[3] ));
 sky130_fd_sc_hd__dfrtp_2 _18785_ (.CLK(clknet_leaf_212_clk),
    .D(_00083_),
    .RESET_B(net274),
    .Q(\center_y[4] ));
 sky130_fd_sc_hd__dfrtp_2 _18786_ (.CLK(clknet_leaf_212_clk),
    .D(_00084_),
    .RESET_B(net274),
    .Q(\center_y[5] ));
 sky130_fd_sc_hd__dfrtp_2 _18787_ (.CLK(clknet_leaf_212_clk),
    .D(_00085_),
    .RESET_B(net274),
    .Q(\center_y[6] ));
 sky130_fd_sc_hd__dfrtp_1 _18788_ (.CLK(clknet_leaf_200_clk),
    .D(_00086_),
    .RESET_B(net270),
    .Q(\shex_center_x[0] ));
 sky130_fd_sc_hd__dfrtp_1 _18789_ (.CLK(clknet_leaf_201_clk),
    .D(_00087_),
    .RESET_B(net271),
    .Q(\shex_center_x[1] ));
 sky130_fd_sc_hd__dfrtp_1 _18790_ (.CLK(clknet_leaf_202_clk),
    .D(_00088_),
    .RESET_B(net276),
    .Q(\shex_center_x[2] ));
 sky130_fd_sc_hd__dfrtp_1 _18791_ (.CLK(clknet_leaf_203_clk),
    .D(_00089_),
    .RESET_B(net277),
    .Q(\shex_center_x[3] ));
 sky130_fd_sc_hd__dfrtp_1 _18792_ (.CLK(clknet_leaf_205_clk),
    .D(_00090_),
    .RESET_B(net276),
    .Q(\shex_center_x[4] ));
 sky130_fd_sc_hd__dfrtp_1 _18793_ (.CLK(clknet_leaf_207_clk),
    .D(_00091_),
    .RESET_B(net278),
    .Q(\shex_center_x[5] ));
 sky130_fd_sc_hd__dfrtp_1 _18794_ (.CLK(clknet_leaf_207_clk),
    .D(_00092_),
    .RESET_B(net278),
    .Q(\shex_center_x[6] ));
 sky130_fd_sc_hd__dfrtp_1 _18795_ (.CLK(clknet_leaf_205_clk),
    .D(_00093_),
    .RESET_B(net277),
    .Q(\shex_center_y[0] ));
 sky130_fd_sc_hd__dfrtp_1 _18796_ (.CLK(clknet_leaf_209_clk),
    .D(_00094_),
    .RESET_B(net273),
    .Q(\shex_center_y[1] ));
 sky130_fd_sc_hd__dfrtp_1 _18797_ (.CLK(clknet_leaf_209_clk),
    .D(_00095_),
    .RESET_B(net273),
    .Q(\shex_center_y[2] ));
 sky130_fd_sc_hd__dfrtp_1 _18798_ (.CLK(clknet_leaf_209_clk),
    .D(_00096_),
    .RESET_B(net275),
    .Q(\shex_center_y[3] ));
 sky130_fd_sc_hd__dfrtp_1 _18799_ (.CLK(clknet_leaf_208_clk),
    .D(_00097_),
    .RESET_B(net278),
    .Q(\shex_center_y[4] ));
 sky130_fd_sc_hd__dfrtp_1 _18800_ (.CLK(clknet_leaf_208_clk),
    .D(_00098_),
    .RESET_B(net278),
    .Q(\shex_center_y[5] ));
 sky130_fd_sc_hd__dfrtp_1 _18801_ (.CLK(clknet_leaf_211_clk),
    .D(_00099_),
    .RESET_B(net275),
    .Q(\shex_center_y[6] ));
 sky130_fd_sc_hd__dfrtp_4 _18802_ (.CLK(clknet_leaf_201_clk),
    .D(_00100_),
    .RESET_B(net270),
    .Q(\cand_x[0] ));
 sky130_fd_sc_hd__dfrtp_4 _18803_ (.CLK(clknet_leaf_199_clk),
    .D(_00101_),
    .RESET_B(net277),
    .Q(\cand_x[1] ));
 sky130_fd_sc_hd__dfrtp_4 _18804_ (.CLK(clknet_leaf_202_clk),
    .D(_00102_),
    .RESET_B(net276),
    .Q(\cand_x[2] ));
 sky130_fd_sc_hd__dfrtp_4 _18805_ (.CLK(clknet_leaf_204_clk),
    .D(_00103_),
    .RESET_B(net277),
    .Q(\cand_x[3] ));
 sky130_fd_sc_hd__dfrtp_4 _18806_ (.CLK(clknet_leaf_204_clk),
    .D(_00104_),
    .RESET_B(net277),
    .Q(\cand_x[4] ));
 sky130_fd_sc_hd__dfrtp_4 _18807_ (.CLK(clknet_leaf_208_clk),
    .D(_00105_),
    .RESET_B(net278),
    .Q(\cand_x[5] ));
 sky130_fd_sc_hd__dfrtp_2 _18808_ (.CLK(clknet_leaf_214_clk),
    .D(_00106_),
    .RESET_B(net274),
    .Q(\cand_x[6] ));
 sky130_fd_sc_hd__dfrtp_4 _18809_ (.CLK(clknet_leaf_205_clk),
    .D(_00107_),
    .RESET_B(net277),
    .Q(\cand_y[0] ));
 sky130_fd_sc_hd__dfrtp_4 _18810_ (.CLK(clknet_leaf_217_clk),
    .D(_00108_),
    .RESET_B(net273),
    .Q(\cand_y[1] ));
 sky130_fd_sc_hd__dfrtp_4 _18811_ (.CLK(clknet_leaf_216_clk),
    .D(_00109_),
    .RESET_B(net273),
    .Q(\cand_y[2] ));
 sky130_fd_sc_hd__dfrtp_4 _18812_ (.CLK(clknet_leaf_216_clk),
    .D(_00110_),
    .RESET_B(net275),
    .Q(\cand_y[3] ));
 sky130_fd_sc_hd__dfrtp_2 _18813_ (.CLK(clknet_5_30__leaf_clk),
    .D(_00111_),
    .RESET_B(net275),
    .Q(\cand_y[4] ));
 sky130_fd_sc_hd__dfrtp_4 _18814_ (.CLK(clknet_leaf_212_clk),
    .D(_00112_),
    .RESET_B(net274),
    .Q(\cand_y[5] ));
 sky130_fd_sc_hd__dfrtp_1 _18815_ (.CLK(clknet_leaf_213_clk),
    .D(_00113_),
    .RESET_B(net274),
    .Q(\cand_y[6] ));
 sky130_fd_sc_hd__dfrtp_1 _18816_ (.CLK(clknet_leaf_226_clk),
    .D(_00114_),
    .RESET_B(net279),
    .Q(\pixel_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _18817_ (.CLK(clknet_leaf_226_clk),
    .D(_00115_),
    .RESET_B(net279),
    .Q(\pixel_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _18818_ (.CLK(clknet_leaf_226_clk),
    .D(_00116_),
    .RESET_B(net279),
    .Q(\pixel_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _18819_ (.CLK(clknet_leaf_226_clk),
    .D(_00117_),
    .RESET_B(net279),
    .Q(\pixel_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _18820_ (.CLK(clknet_leaf_225_clk),
    .D(_00118_),
    .RESET_B(net279),
    .Q(\pixel_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _18821_ (.CLK(clknet_leaf_223_clk),
    .D(_00119_),
    .RESET_B(net279),
    .Q(\pixel_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _18822_ (.CLK(clknet_leaf_221_clk),
    .D(_00120_),
    .RESET_B(net279),
    .Q(\pixel_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _18823_ (.CLK(clknet_leaf_225_clk),
    .D(_00121_),
    .RESET_B(net279),
    .Q(\pixel_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _18824_ (.CLK(clknet_leaf_197_clk),
    .D(_00122_),
    .RESET_B(net266),
    .Q(\pixel_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_2 _18825_ (.CLK(clknet_leaf_200_clk),
    .D(_00123_),
    .RESET_B(net270),
    .Q(\point_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _18826_ (.CLK(clknet_leaf_200_clk),
    .D(_00124_),
    .RESET_B(net270),
    .Q(\point_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _18827_ (.CLK(clknet_leaf_199_clk),
    .D(_00125_),
    .RESET_B(net277),
    .Q(\point_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _18828_ (.CLK(clknet_leaf_199_clk),
    .D(_00126_),
    .RESET_B(net270),
    .Q(\point_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_2 _18829_ (.CLK(clknet_leaf_198_clk),
    .D(_00127_),
    .RESET_B(net267),
    .Q(shex_load));
 sky130_fd_sc_hd__dfxtp_1 _18830_ (.CLK(clknet_leaf_185_clk),
    .D(_00128_),
    .Q(\current_accum_sad[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18831_ (.CLK(clknet_leaf_186_clk),
    .D(_00129_),
    .Q(\current_accum_sad[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18832_ (.CLK(clknet_leaf_186_clk),
    .D(_00130_),
    .Q(\current_accum_sad[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18833_ (.CLK(clknet_leaf_187_clk),
    .D(_00131_),
    .Q(\current_accum_sad[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18834_ (.CLK(clknet_leaf_187_clk),
    .D(_00132_),
    .Q(\current_accum_sad[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18835_ (.CLK(clknet_leaf_187_clk),
    .D(_00133_),
    .Q(\current_accum_sad[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18836_ (.CLK(clknet_leaf_186_clk),
    .D(_00134_),
    .Q(\current_accum_sad[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18837_ (.CLK(clknet_leaf_191_clk),
    .D(_00135_),
    .Q(\current_accum_sad[7] ));
 sky130_fd_sc_hd__dfxtp_1 _18838_ (.CLK(clknet_leaf_189_clk),
    .D(_00136_),
    .Q(\current_accum_sad[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18839_ (.CLK(clknet_leaf_189_clk),
    .D(_00137_),
    .Q(\current_accum_sad[9] ));
 sky130_fd_sc_hd__dfxtp_1 _18840_ (.CLK(clknet_leaf_200_clk),
    .D(_00138_),
    .Q(\current_accum_sad[10] ));
 sky130_fd_sc_hd__dfxtp_1 _18841_ (.CLK(clknet_leaf_200_clk),
    .D(_00139_),
    .Q(\current_accum_sad[11] ));
 sky130_fd_sc_hd__dfxtp_1 _18842_ (.CLK(clknet_leaf_200_clk),
    .D(_00140_),
    .Q(\current_accum_sad[12] ));
 sky130_fd_sc_hd__dfxtp_1 _18843_ (.CLK(clknet_leaf_194_clk),
    .D(_00141_),
    .Q(\current_accum_sad[13] ));
 sky130_fd_sc_hd__dfxtp_1 _18844_ (.CLK(clknet_leaf_194_clk),
    .D(_00142_),
    .Q(\current_accum_sad[14] ));
 sky130_fd_sc_hd__dfxtp_1 _18845_ (.CLK(clknet_leaf_198_clk),
    .D(_00143_),
    .Q(\current_accum_sad[15] ));
 sky130_fd_sc_hd__dfxtp_1 _18846_ (.CLK(clknet_leaf_205_clk),
    .D(_00144_),
    .Q(\best_cand_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18847_ (.CLK(clknet_leaf_214_clk),
    .D(_00145_),
    .Q(\best_cand_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18848_ (.CLK(clknet_leaf_216_clk),
    .D(_00146_),
    .Q(\best_cand_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18849_ (.CLK(clknet_leaf_214_clk),
    .D(_00147_),
    .Q(\best_cand_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18850_ (.CLK(clknet_leaf_212_clk),
    .D(_00148_),
    .Q(\best_cand_y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18851_ (.CLK(clknet_leaf_213_clk),
    .D(_00149_),
    .Q(\best_cand_y[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18852_ (.CLK(clknet_leaf_213_clk),
    .D(_00150_),
    .Q(\best_cand_y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18853_ (.CLK(clknet_leaf_180_clk),
    .D(_00151_),
    .Q(\cur_mb_mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18854_ (.CLK(clknet_leaf_181_clk),
    .D(_00152_),
    .Q(\cur_mb_mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18855_ (.CLK(clknet_leaf_184_clk),
    .D(_00153_),
    .Q(\cur_mb_mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18856_ (.CLK(clknet_leaf_180_clk),
    .D(_00154_),
    .Q(\cur_mb_mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18857_ (.CLK(clknet_leaf_183_clk),
    .D(_00155_),
    .Q(\cur_mb_mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18858_ (.CLK(clknet_leaf_183_clk),
    .D(_00156_),
    .Q(\cur_mb_mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18859_ (.CLK(clknet_leaf_180_clk),
    .D(_00157_),
    .Q(\cur_mb_mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18860_ (.CLK(clknet_leaf_184_clk),
    .D(_00158_),
    .Q(\cur_mb_mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18861_ (.CLK(clknet_leaf_98_clk),
    .D(_00159_),
    .Q(\cur_mb_mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _18862_ (.CLK(clknet_leaf_116_clk),
    .D(_00160_),
    .Q(\cur_mb_mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18863_ (.CLK(clknet_leaf_104_clk),
    .D(_00161_),
    .Q(\cur_mb_mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18864_ (.CLK(clknet_leaf_102_clk),
    .D(_00162_),
    .Q(\cur_mb_mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18865_ (.CLK(clknet_leaf_120_clk),
    .D(_00163_),
    .Q(\cur_mb_mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18866_ (.CLK(clknet_leaf_183_clk),
    .D(_00164_),
    .Q(\cur_mb_mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18867_ (.CLK(clknet_leaf_177_clk),
    .D(_00165_),
    .Q(\cur_mb_mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _18868_ (.CLK(clknet_leaf_177_clk),
    .D(_00166_),
    .Q(\cur_mb_mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18869_ (.CLK(clknet_leaf_101_clk),
    .D(_00167_),
    .Q(\cur_mb_mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18870_ (.CLK(clknet_leaf_104_clk),
    .D(_00168_),
    .Q(\cur_mb_mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18871_ (.CLK(clknet_leaf_100_clk),
    .D(_00169_),
    .Q(\cur_mb_mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18872_ (.CLK(clknet_leaf_99_clk),
    .D(_00170_),
    .Q(\cur_mb_mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18873_ (.CLK(clknet_leaf_121_clk),
    .D(_00171_),
    .Q(\cur_mb_mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18874_ (.CLK(clknet_leaf_117_clk),
    .D(_00172_),
    .Q(\cur_mb_mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18875_ (.CLK(clknet_leaf_177_clk),
    .D(_00173_),
    .Q(\cur_mb_mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _18876_ (.CLK(clknet_leaf_184_clk),
    .D(_00174_),
    .Q(\cur_mb_mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18877_ (.CLK(clknet_leaf_44_clk),
    .D(_00175_),
    .Q(\cur_mb_mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18878_ (.CLK(clknet_leaf_61_clk),
    .D(_00176_),
    .Q(\cur_mb_mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18879_ (.CLK(clknet_leaf_51_clk),
    .D(_00177_),
    .Q(\cur_mb_mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18880_ (.CLK(clknet_leaf_44_clk),
    .D(_00178_),
    .Q(\cur_mb_mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18881_ (.CLK(clknet_leaf_121_clk),
    .D(_00179_),
    .Q(\cur_mb_mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18882_ (.CLK(clknet_leaf_122_clk),
    .D(_00180_),
    .Q(\cur_mb_mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18883_ (.CLK(clknet_leaf_147_clk),
    .D(_00181_),
    .Q(\cur_mb_mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18884_ (.CLK(clknet_leaf_184_clk),
    .D(_00182_),
    .Q(\cur_mb_mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18885_ (.CLK(clknet_leaf_111_clk),
    .D(_00183_),
    .Q(\cur_mb_mem[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18886_ (.CLK(clknet_leaf_123_clk),
    .D(_00184_),
    .Q(\cur_mb_mem[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18887_ (.CLK(clknet_leaf_120_clk),
    .D(_00185_),
    .Q(\cur_mb_mem[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18888_ (.CLK(clknet_leaf_116_clk),
    .D(_00186_),
    .Q(\cur_mb_mem[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18889_ (.CLK(clknet_leaf_183_clk),
    .D(_00187_),
    .Q(\cur_mb_mem[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18890_ (.CLK(clknet_leaf_183_clk),
    .D(_00188_),
    .Q(\cur_mb_mem[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _18891_ (.CLK(clknet_leaf_178_clk),
    .D(_00189_),
    .Q(\cur_mb_mem[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18892_ (.CLK(clknet_leaf_183_clk),
    .D(_00190_),
    .Q(\cur_mb_mem[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18893_ (.CLK(clknet_leaf_100_clk),
    .D(_00191_),
    .Q(\cur_mb_mem[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18894_ (.CLK(clknet_leaf_115_clk),
    .D(_00192_),
    .Q(\cur_mb_mem[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18895_ (.CLK(clknet_leaf_100_clk),
    .D(_00193_),
    .Q(\cur_mb_mem[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18896_ (.CLK(clknet_leaf_99_clk),
    .D(_00194_),
    .Q(\cur_mb_mem[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18897_ (.CLK(clknet_leaf_178_clk),
    .D(_00195_),
    .Q(\cur_mb_mem[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18898_ (.CLK(clknet_leaf_182_clk),
    .D(_00196_),
    .Q(\cur_mb_mem[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18899_ (.CLK(clknet_leaf_325_clk),
    .D(_00197_),
    .Q(\cur_mb_mem[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18900_ (.CLK(clknet_leaf_325_clk),
    .D(_00198_),
    .Q(\cur_mb_mem[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18901_ (.CLK(clknet_leaf_1_clk),
    .D(_00199_),
    .Q(\cur_mb_mem[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18902_ (.CLK(clknet_leaf_348_clk),
    .D(_00200_),
    .Q(\cur_mb_mem[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18903_ (.CLK(clknet_leaf_1_clk),
    .D(_00201_),
    .Q(\cur_mb_mem[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18904_ (.CLK(clknet_leaf_1_clk),
    .D(_00202_),
    .Q(\cur_mb_mem[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18905_ (.CLK(clknet_leaf_45_clk),
    .D(_00203_),
    .Q(\cur_mb_mem[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18906_ (.CLK(clknet_leaf_44_clk),
    .D(_00204_),
    .Q(\cur_mb_mem[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18907_ (.CLK(clknet_leaf_49_clk),
    .D(_00205_),
    .Q(\cur_mb_mem[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18908_ (.CLK(clknet_leaf_325_clk),
    .D(_00206_),
    .Q(\cur_mb_mem[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18909_ (.CLK(clknet_leaf_313_clk),
    .D(_00207_),
    .Q(\cur_mb_mem[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18910_ (.CLK(clknet_leaf_254_clk),
    .D(_00208_),
    .Q(\cur_mb_mem[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18911_ (.CLK(clknet_leaf_314_clk),
    .D(_00209_),
    .Q(\cur_mb_mem[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18912_ (.CLK(clknet_leaf_249_clk),
    .D(_00210_),
    .Q(\cur_mb_mem[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18913_ (.CLK(clknet_leaf_181_clk),
    .D(_00211_),
    .Q(\cur_mb_mem[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18914_ (.CLK(clknet_leaf_181_clk),
    .D(_00212_),
    .Q(\cur_mb_mem[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18915_ (.CLK(clknet_leaf_321_clk),
    .D(_00213_),
    .Q(\cur_mb_mem[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18916_ (.CLK(clknet_leaf_321_clk),
    .D(_00214_),
    .Q(\cur_mb_mem[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18917_ (.CLK(clknet_leaf_1_clk),
    .D(_00215_),
    .Q(\cur_mb_mem[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18918_ (.CLK(clknet_leaf_335_clk),
    .D(_00216_),
    .Q(\cur_mb_mem[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18919_ (.CLK(clknet_leaf_1_clk),
    .D(_00217_),
    .Q(\cur_mb_mem[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18920_ (.CLK(clknet_leaf_9_clk),
    .D(_00218_),
    .Q(\cur_mb_mem[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18921_ (.CLK(clknet_leaf_120_clk),
    .D(_00219_),
    .Q(\cur_mb_mem[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18922_ (.CLK(clknet_leaf_117_clk),
    .D(_00220_),
    .Q(\cur_mb_mem[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18923_ (.CLK(clknet_leaf_336_clk),
    .D(_00221_),
    .Q(\cur_mb_mem[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18924_ (.CLK(clknet_leaf_330_clk),
    .D(_00222_),
    .Q(\cur_mb_mem[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18925_ (.CLK(clknet_leaf_8_clk),
    .D(_00223_),
    .Q(\cur_mb_mem[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18926_ (.CLK(clknet_leaf_345_clk),
    .D(_00224_),
    .Q(\cur_mb_mem[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18927_ (.CLK(clknet_leaf_11_clk),
    .D(_00225_),
    .Q(\cur_mb_mem[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18928_ (.CLK(clknet_leaf_8_clk),
    .D(_00226_),
    .Q(\cur_mb_mem[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18929_ (.CLK(clknet_leaf_120_clk),
    .D(_00227_),
    .Q(\cur_mb_mem[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18930_ (.CLK(clknet_leaf_116_clk),
    .D(_00228_),
    .Q(\cur_mb_mem[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18931_ (.CLK(clknet_leaf_338_clk),
    .D(_00229_),
    .Q(\cur_mb_mem[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18932_ (.CLK(clknet_leaf_324_clk),
    .D(_00230_),
    .Q(\cur_mb_mem[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18933_ (.CLK(clknet_leaf_3_clk),
    .D(_00231_),
    .Q(\cur_mb_mem[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18934_ (.CLK(clknet_leaf_379_clk),
    .D(_00232_),
    .Q(\cur_mb_mem[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18935_ (.CLK(clknet_leaf_2_clk),
    .D(_00233_),
    .Q(\cur_mb_mem[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18936_ (.CLK(clknet_leaf_3_clk),
    .D(_00234_),
    .Q(\cur_mb_mem[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18937_ (.CLK(clknet_leaf_355_clk),
    .D(_00235_),
    .Q(\cur_mb_mem[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18938_ (.CLK(clknet_leaf_350_clk),
    .D(_00236_),
    .Q(\cur_mb_mem[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18939_ (.CLK(clknet_leaf_154_clk),
    .D(_00237_),
    .Q(\cur_mb_mem[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18940_ (.CLK(clknet_leaf_337_clk),
    .D(_00238_),
    .Q(\cur_mb_mem[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18941_ (.CLK(clknet_leaf_243_clk),
    .D(_00239_),
    .Q(\cur_mb_mem[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18942_ (.CLK(clknet_leaf_47_clk),
    .D(_00240_),
    .Q(\cur_mb_mem[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18943_ (.CLK(clknet_leaf_244_clk),
    .D(_00241_),
    .Q(\cur_mb_mem[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18944_ (.CLK(clknet_leaf_246_clk),
    .D(_00242_),
    .Q(\cur_mb_mem[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18945_ (.CLK(clknet_leaf_237_clk),
    .D(_00243_),
    .Q(\cur_mb_mem[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18946_ (.CLK(clknet_leaf_156_clk),
    .D(_00244_),
    .Q(\cur_mb_mem[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18947_ (.CLK(clknet_leaf_334_clk),
    .D(_00245_),
    .Q(\cur_mb_mem[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18948_ (.CLK(clknet_leaf_156_clk),
    .D(_00246_),
    .Q(\cur_mb_mem[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18949_ (.CLK(clknet_leaf_175_clk),
    .D(_00247_),
    .Q(\cur_mb_mem[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18950_ (.CLK(clknet_leaf_149_clk),
    .D(_00248_),
    .Q(\cur_mb_mem[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18951_ (.CLK(clknet_leaf_175_clk),
    .D(_00249_),
    .Q(\cur_mb_mem[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18952_ (.CLK(clknet_leaf_175_clk),
    .D(_00250_),
    .Q(\cur_mb_mem[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18953_ (.CLK(clknet_leaf_181_clk),
    .D(_00251_),
    .Q(\cur_mb_mem[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18954_ (.CLK(clknet_leaf_182_clk),
    .D(_00252_),
    .Q(\cur_mb_mem[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18955_ (.CLK(clknet_leaf_149_clk),
    .D(_00253_),
    .Q(\cur_mb_mem[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18956_ (.CLK(clknet_leaf_159_clk),
    .D(_00254_),
    .Q(\cur_mb_mem[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18957_ (.CLK(clknet_leaf_46_clk),
    .D(_00255_),
    .Q(\cur_mb_mem[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18958_ (.CLK(clknet_leaf_338_clk),
    .D(_00256_),
    .Q(\cur_mb_mem[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18959_ (.CLK(clknet_leaf_46_clk),
    .D(_00257_),
    .Q(\cur_mb_mem[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18960_ (.CLK(clknet_leaf_46_clk),
    .D(_00258_),
    .Q(\cur_mb_mem[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18961_ (.CLK(clknet_leaf_331_clk),
    .D(_00259_),
    .Q(\cur_mb_mem[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18962_ (.CLK(clknet_leaf_331_clk),
    .D(_00260_),
    .Q(\cur_mb_mem[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18963_ (.CLK(clknet_leaf_323_clk),
    .D(_00261_),
    .Q(\cur_mb_mem[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18964_ (.CLK(clknet_leaf_242_clk),
    .D(_00262_),
    .Q(\cur_mb_mem[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18965_ (.CLK(clknet_leaf_353_clk),
    .D(_00263_),
    .Q(\cur_mb_mem[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18966_ (.CLK(clknet_leaf_52_clk),
    .D(_00264_),
    .Q(\cur_mb_mem[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18967_ (.CLK(clknet_leaf_353_clk),
    .D(_00265_),
    .Q(\cur_mb_mem[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18968_ (.CLK(clknet_leaf_353_clk),
    .D(_00266_),
    .Q(\cur_mb_mem[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18969_ (.CLK(clknet_leaf_124_clk),
    .D(_00267_),
    .Q(\cur_mb_mem[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18970_ (.CLK(clknet_leaf_119_clk),
    .D(_00268_),
    .Q(\cur_mb_mem[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18971_ (.CLK(clknet_leaf_335_clk),
    .D(_00269_),
    .Q(\cur_mb_mem[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18972_ (.CLK(clknet_leaf_176_clk),
    .D(_00270_),
    .Q(\cur_mb_mem[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18973_ (.CLK(clknet_leaf_253_clk),
    .D(_00271_),
    .Q(\cur_mb_mem[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18974_ (.CLK(clknet_leaf_252_clk),
    .D(_00272_),
    .Q(\cur_mb_mem[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18975_ (.CLK(clknet_leaf_261_clk),
    .D(_00273_),
    .Q(\cur_mb_mem[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18976_ (.CLK(clknet_leaf_253_clk),
    .D(_00274_),
    .Q(\cur_mb_mem[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _18977_ (.CLK(clknet_leaf_148_clk),
    .D(_00275_),
    .Q(\cur_mb_mem[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18978_ (.CLK(clknet_leaf_148_clk),
    .D(_00276_),
    .Q(\cur_mb_mem[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18979_ (.CLK(clknet_leaf_149_clk),
    .D(_00277_),
    .Q(\cur_mb_mem[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18980_ (.CLK(clknet_leaf_156_clk),
    .D(_00278_),
    .Q(\cur_mb_mem[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18981_ (.CLK(clknet_leaf_245_clk),
    .D(_00279_),
    .Q(\cur_mb_mem[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18982_ (.CLK(clknet_leaf_53_clk),
    .D(_00280_),
    .Q(\cur_mb_mem[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18983_ (.CLK(clknet_leaf_244_clk),
    .D(_00281_),
    .Q(\cur_mb_mem[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18984_ (.CLK(clknet_leaf_246_clk),
    .D(_00282_),
    .Q(\cur_mb_mem[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18985_ (.CLK(clknet_leaf_180_clk),
    .D(_00283_),
    .Q(\cur_mb_mem[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18986_ (.CLK(clknet_leaf_182_clk),
    .D(_00284_),
    .Q(\cur_mb_mem[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18987_ (.CLK(clknet_leaf_49_clk),
    .D(_00285_),
    .Q(\cur_mb_mem[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18988_ (.CLK(clknet_leaf_47_clk),
    .D(_00286_),
    .Q(\cur_mb_mem[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18989_ (.CLK(clknet_leaf_173_clk),
    .D(_00287_),
    .Q(\cur_mb_mem[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18990_ (.CLK(clknet_leaf_241_clk),
    .D(_00288_),
    .Q(\cur_mb_mem[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18991_ (.CLK(clknet_leaf_173_clk),
    .D(_00289_),
    .Q(\cur_mb_mem[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18992_ (.CLK(clknet_leaf_123_clk),
    .D(_00290_),
    .Q(\cur_mb_mem[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18993_ (.CLK(clknet_leaf_181_clk),
    .D(_00291_),
    .Q(\cur_mb_mem[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18994_ (.CLK(clknet_leaf_182_clk),
    .D(_00292_),
    .Q(\cur_mb_mem[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18995_ (.CLK(clknet_leaf_239_clk),
    .D(_00293_),
    .Q(\cur_mb_mem[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18996_ (.CLK(clknet_leaf_238_clk),
    .D(_00294_),
    .Q(\cur_mb_mem[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18997_ (.CLK(clknet_leaf_97_clk),
    .D(_00295_),
    .Q(\cur_mb_mem[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18998_ (.CLK(clknet_leaf_233_clk),
    .D(_00296_),
    .Q(\cur_mb_mem[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18999_ (.CLK(clknet_leaf_97_clk),
    .D(_00297_),
    .Q(\cur_mb_mem[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19000_ (.CLK(clknet_leaf_104_clk),
    .D(_00298_),
    .Q(\cur_mb_mem[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19001_ (.CLK(clknet_leaf_181_clk),
    .D(_00299_),
    .Q(\cur_mb_mem[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19002_ (.CLK(clknet_leaf_182_clk),
    .D(_00300_),
    .Q(\cur_mb_mem[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19003_ (.CLK(clknet_leaf_154_clk),
    .D(_00301_),
    .Q(\cur_mb_mem[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19004_ (.CLK(clknet_leaf_141_clk),
    .D(_00302_),
    .Q(\cur_mb_mem[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19005_ (.CLK(clknet_leaf_109_clk),
    .D(_00303_),
    .Q(\cur_mb_mem[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19006_ (.CLK(clknet_leaf_38_clk),
    .D(_00304_),
    .Q(\cur_mb_mem[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19007_ (.CLK(clknet_leaf_131_clk),
    .D(_00305_),
    .Q(\cur_mb_mem[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19008_ (.CLK(clknet_leaf_115_clk),
    .D(_00306_),
    .Q(\cur_mb_mem[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19009_ (.CLK(clknet_leaf_120_clk),
    .D(_00307_),
    .Q(\cur_mb_mem[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19010_ (.CLK(clknet_leaf_123_clk),
    .D(_00308_),
    .Q(\cur_mb_mem[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19011_ (.CLK(clknet_leaf_337_clk),
    .D(_00309_),
    .Q(\cur_mb_mem[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19012_ (.CLK(clknet_leaf_149_clk),
    .D(_00310_),
    .Q(\cur_mb_mem[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19013_ (.CLK(clknet_leaf_174_clk),
    .D(_00311_),
    .Q(\cur_mb_mem[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19014_ (.CLK(clknet_leaf_238_clk),
    .D(_00312_),
    .Q(\cur_mb_mem[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19015_ (.CLK(clknet_leaf_174_clk),
    .D(_00313_),
    .Q(\cur_mb_mem[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19016_ (.CLK(clknet_leaf_170_clk),
    .D(_00314_),
    .Q(\cur_mb_mem[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19017_ (.CLK(clknet_leaf_237_clk),
    .D(_00315_),
    .Q(\cur_mb_mem[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19018_ (.CLK(clknet_leaf_156_clk),
    .D(_00316_),
    .Q(\cur_mb_mem[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19019_ (.CLK(clknet_leaf_238_clk),
    .D(_00317_),
    .Q(\cur_mb_mem[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19020_ (.CLK(clknet_leaf_161_clk),
    .D(_00318_),
    .Q(\cur_mb_mem[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19021_ (.CLK(clknet_leaf_34_clk),
    .D(_00319_),
    .Q(\cur_mb_mem[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19022_ (.CLK(clknet_leaf_39_clk),
    .D(_00320_),
    .Q(\cur_mb_mem[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19023_ (.CLK(clknet_leaf_27_clk),
    .D(_00321_),
    .Q(\cur_mb_mem[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19024_ (.CLK(clknet_leaf_27_clk),
    .D(_00322_),
    .Q(\cur_mb_mem[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19025_ (.CLK(clknet_leaf_332_clk),
    .D(_00323_),
    .Q(\cur_mb_mem[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19026_ (.CLK(clknet_leaf_332_clk),
    .D(_00324_),
    .Q(\cur_mb_mem[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19027_ (.CLK(clknet_leaf_48_clk),
    .D(_00325_),
    .Q(\cur_mb_mem[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19028_ (.CLK(clknet_leaf_343_clk),
    .D(_00326_),
    .Q(\cur_mb_mem[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19029_ (.CLK(clknet_leaf_170_clk),
    .D(_00327_),
    .Q(\cur_mb_mem[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19030_ (.CLK(clknet_leaf_338_clk),
    .D(_00328_),
    .Q(\cur_mb_mem[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19031_ (.CLK(clknet_leaf_166_clk),
    .D(_00329_),
    .Q(\cur_mb_mem[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19032_ (.CLK(clknet_leaf_170_clk),
    .D(_00330_),
    .Q(\cur_mb_mem[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19033_ (.CLK(clknet_leaf_123_clk),
    .D(_00331_),
    .Q(\cur_mb_mem[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19034_ (.CLK(clknet_leaf_124_clk),
    .D(_00332_),
    .Q(\cur_mb_mem[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19035_ (.CLK(clknet_leaf_340_clk),
    .D(_00333_),
    .Q(\cur_mb_mem[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19036_ (.CLK(clknet_leaf_145_clk),
    .D(_00334_),
    .Q(\cur_mb_mem[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19037_ (.CLK(clknet_leaf_252_clk),
    .D(_00335_),
    .Q(\cur_mb_mem[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19038_ (.CLK(clknet_leaf_233_clk),
    .D(_00336_),
    .Q(\cur_mb_mem[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19039_ (.CLK(clknet_leaf_234_clk),
    .D(_00337_),
    .Q(\cur_mb_mem[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19040_ (.CLK(clknet_leaf_193_clk),
    .D(_00338_),
    .Q(\cur_mb_mem[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19041_ (.CLK(clknet_leaf_180_clk),
    .D(_00339_),
    .Q(\cur_mb_mem[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19042_ (.CLK(clknet_leaf_179_clk),
    .D(_00340_),
    .Q(\cur_mb_mem[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19043_ (.CLK(clknet_leaf_320_clk),
    .D(_00341_),
    .Q(\cur_mb_mem[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19044_ (.CLK(clknet_leaf_320_clk),
    .D(_00342_),
    .Q(\cur_mb_mem[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19045_ (.CLK(clknet_leaf_173_clk),
    .D(_00343_),
    .Q(\cur_mb_mem[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19046_ (.CLK(clknet_leaf_126_clk),
    .D(_00344_),
    .Q(\cur_mb_mem[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19047_ (.CLK(clknet_leaf_173_clk),
    .D(_00345_),
    .Q(\cur_mb_mem[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19048_ (.CLK(clknet_leaf_123_clk),
    .D(_00346_),
    .Q(\cur_mb_mem[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19049_ (.CLK(clknet_leaf_122_clk),
    .D(_00347_),
    .Q(\cur_mb_mem[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19050_ (.CLK(clknet_leaf_122_clk),
    .D(_00348_),
    .Q(\cur_mb_mem[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19051_ (.CLK(clknet_leaf_128_clk),
    .D(_00349_),
    .Q(\cur_mb_mem[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19052_ (.CLK(clknet_leaf_128_clk),
    .D(_00350_),
    .Q(\cur_mb_mem[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19053_ (.CLK(clknet_leaf_172_clk),
    .D(_00351_),
    .Q(\cur_mb_mem[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19054_ (.CLK(clknet_leaf_172_clk),
    .D(_00352_),
    .Q(\cur_mb_mem[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19055_ (.CLK(clknet_leaf_172_clk),
    .D(_00353_),
    .Q(\cur_mb_mem[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19056_ (.CLK(clknet_leaf_185_clk),
    .D(_00354_),
    .Q(\cur_mb_mem[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19057_ (.CLK(clknet_leaf_121_clk),
    .D(_00355_),
    .Q(\cur_mb_mem[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19058_ (.CLK(clknet_leaf_117_clk),
    .D(_00356_),
    .Q(\cur_mb_mem[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19059_ (.CLK(clknet_leaf_177_clk),
    .D(_00357_),
    .Q(\cur_mb_mem[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19060_ (.CLK(clknet_leaf_125_clk),
    .D(_00358_),
    .Q(\cur_mb_mem[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19061_ (.CLK(clknet_leaf_179_clk),
    .D(_00359_),
    .Q(\cur_mb_mem[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19062_ (.CLK(clknet_leaf_177_clk),
    .D(_00360_),
    .Q(\cur_mb_mem[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19063_ (.CLK(clknet_leaf_171_clk),
    .D(_00361_),
    .Q(\cur_mb_mem[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19064_ (.CLK(clknet_leaf_171_clk),
    .D(_00362_),
    .Q(\cur_mb_mem[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19065_ (.CLK(clknet_leaf_122_clk),
    .D(_00363_),
    .Q(\cur_mb_mem[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19066_ (.CLK(clknet_leaf_122_clk),
    .D(_00364_),
    .Q(\cur_mb_mem[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19067_ (.CLK(clknet_leaf_128_clk),
    .D(_00365_),
    .Q(\cur_mb_mem[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19068_ (.CLK(clknet_leaf_126_clk),
    .D(_00366_),
    .Q(\cur_mb_mem[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19069_ (.CLK(clknet_leaf_109_clk),
    .D(_00367_),
    .Q(\cur_mb_mem[27][0] ));
 sky130_fd_sc_hd__dfxtp_2 _19070_ (.CLK(clknet_leaf_135_clk),
    .D(_00368_),
    .Q(\cur_mb_mem[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19071_ (.CLK(clknet_leaf_135_clk),
    .D(_00369_),
    .Q(\cur_mb_mem[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19072_ (.CLK(clknet_leaf_116_clk),
    .D(_00370_),
    .Q(\cur_mb_mem[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19073_ (.CLK(clknet_leaf_121_clk),
    .D(_00371_),
    .Q(\cur_mb_mem[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19074_ (.CLK(clknet_leaf_122_clk),
    .D(_00372_),
    .Q(\cur_mb_mem[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19075_ (.CLK(clknet_leaf_129_clk),
    .D(_00373_),
    .Q(\cur_mb_mem[27][6] ));
 sky130_fd_sc_hd__dfxtp_4 _19076_ (.CLK(clknet_leaf_125_clk),
    .D(_00374_),
    .Q(\cur_mb_mem[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19077_ (.CLK(clknet_leaf_173_clk),
    .D(_00375_),
    .Q(\cur_mb_mem[28][0] ));
 sky130_fd_sc_hd__dfxtp_2 _19078_ (.CLK(clknet_leaf_172_clk),
    .D(_00376_),
    .Q(\cur_mb_mem[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19079_ (.CLK(clknet_leaf_173_clk),
    .D(_00377_),
    .Q(\cur_mb_mem[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19080_ (.CLK(clknet_leaf_185_clk),
    .D(_00378_),
    .Q(\cur_mb_mem[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19081_ (.CLK(clknet_leaf_123_clk),
    .D(_00379_),
    .Q(\cur_mb_mem[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19082_ (.CLK(clknet_leaf_123_clk),
    .D(_00380_),
    .Q(\cur_mb_mem[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19083_ (.CLK(clknet_leaf_128_clk),
    .D(_00381_),
    .Q(\cur_mb_mem[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19084_ (.CLK(clknet_leaf_180_clk),
    .D(_00382_),
    .Q(\cur_mb_mem[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19085_ (.CLK(clknet_leaf_110_clk),
    .D(_00383_),
    .Q(\cur_mb_mem[29][0] ));
 sky130_fd_sc_hd__dfxtp_2 _19086_ (.CLK(clknet_leaf_177_clk),
    .D(_00384_),
    .Q(\cur_mb_mem[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19087_ (.CLK(clknet_leaf_131_clk),
    .D(_00385_),
    .Q(\cur_mb_mem[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19088_ (.CLK(clknet_leaf_116_clk),
    .D(_00386_),
    .Q(\cur_mb_mem[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19089_ (.CLK(clknet_leaf_121_clk),
    .D(_00387_),
    .Q(\cur_mb_mem[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19090_ (.CLK(clknet_leaf_122_clk),
    .D(_00388_),
    .Q(\cur_mb_mem[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19091_ (.CLK(clknet_leaf_128_clk),
    .D(_00389_),
    .Q(\cur_mb_mem[29][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19092_ (.CLK(clknet_leaf_119_clk),
    .D(_00390_),
    .Q(\cur_mb_mem[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19093_ (.CLK(clknet_leaf_100_clk),
    .D(_00391_),
    .Q(\cur_mb_mem[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19094_ (.CLK(clknet_leaf_126_clk),
    .D(_00392_),
    .Q(\cur_mb_mem[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19095_ (.CLK(clknet_leaf_100_clk),
    .D(_00393_),
    .Q(\cur_mb_mem[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19096_ (.CLK(clknet_leaf_99_clk),
    .D(_00394_),
    .Q(\cur_mb_mem[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19097_ (.CLK(clknet_leaf_122_clk),
    .D(_00395_),
    .Q(\cur_mb_mem[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19098_ (.CLK(clknet_leaf_122_clk),
    .D(_00396_),
    .Q(\cur_mb_mem[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19099_ (.CLK(clknet_leaf_128_clk),
    .D(_00397_),
    .Q(\cur_mb_mem[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19100_ (.CLK(clknet_leaf_114_clk),
    .D(_00398_),
    .Q(\cur_mb_mem[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19101_ (.CLK(clknet_leaf_174_clk),
    .D(_00399_),
    .Q(\cur_mb_mem[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19102_ (.CLK(clknet_leaf_175_clk),
    .D(_00400_),
    .Q(\cur_mb_mem[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19103_ (.CLK(clknet_leaf_170_clk),
    .D(_00401_),
    .Q(\cur_mb_mem[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19104_ (.CLK(clknet_leaf_170_clk),
    .D(_00402_),
    .Q(\cur_mb_mem[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19105_ (.CLK(clknet_leaf_135_clk),
    .D(_00403_),
    .Q(\cur_mb_mem[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19106_ (.CLK(clknet_leaf_135_clk),
    .D(_00404_),
    .Q(\cur_mb_mem[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19107_ (.CLK(clknet_leaf_175_clk),
    .D(_00405_),
    .Q(\cur_mb_mem[31][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19108_ (.CLK(clknet_leaf_173_clk),
    .D(_00406_),
    .Q(\cur_mb_mem[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19109_ (.CLK(clknet_leaf_96_clk),
    .D(_00407_),
    .Q(\cur_mb_mem[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19110_ (.CLK(clknet_leaf_136_clk),
    .D(_00408_),
    .Q(\cur_mb_mem[32][1] ));
 sky130_fd_sc_hd__dfxtp_2 _19111_ (.CLK(clknet_leaf_97_clk),
    .D(_00409_),
    .Q(\cur_mb_mem[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19112_ (.CLK(clknet_leaf_97_clk),
    .D(_00410_),
    .Q(\cur_mb_mem[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19113_ (.CLK(clknet_leaf_109_clk),
    .D(_00411_),
    .Q(\cur_mb_mem[32][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19114_ (.CLK(clknet_leaf_109_clk),
    .D(_00412_),
    .Q(\cur_mb_mem[32][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19115_ (.CLK(clknet_leaf_129_clk),
    .D(_00413_),
    .Q(\cur_mb_mem[32][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19116_ (.CLK(clknet_leaf_128_clk),
    .D(_00414_),
    .Q(\cur_mb_mem[32][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19117_ (.CLK(clknet_leaf_95_clk),
    .D(_00415_),
    .Q(\cur_mb_mem[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19118_ (.CLK(clknet_leaf_136_clk),
    .D(_00416_),
    .Q(\cur_mb_mem[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19119_ (.CLK(clknet_leaf_95_clk),
    .D(_00417_),
    .Q(\cur_mb_mem[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19120_ (.CLK(clknet_leaf_96_clk),
    .D(_00418_),
    .Q(\cur_mb_mem[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19121_ (.CLK(clknet_leaf_136_clk),
    .D(_00419_),
    .Q(\cur_mb_mem[33][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19122_ (.CLK(clknet_leaf_136_clk),
    .D(_00420_),
    .Q(\cur_mb_mem[33][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19123_ (.CLK(clknet_leaf_176_clk),
    .D(_00421_),
    .Q(\cur_mb_mem[33][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19124_ (.CLK(clknet_leaf_177_clk),
    .D(_00422_),
    .Q(\cur_mb_mem[33][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19125_ (.CLK(clknet_leaf_245_clk),
    .D(_00423_),
    .Q(\cur_mb_mem[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19126_ (.CLK(clknet_leaf_330_clk),
    .D(_00424_),
    .Q(\cur_mb_mem[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19127_ (.CLK(clknet_leaf_43_clk),
    .D(_00425_),
    .Q(\cur_mb_mem[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19128_ (.CLK(clknet_leaf_246_clk),
    .D(_00426_),
    .Q(\cur_mb_mem[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19129_ (.CLK(clknet_leaf_44_clk),
    .D(_00427_),
    .Q(\cur_mb_mem[34][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19130_ (.CLK(clknet_leaf_57_clk),
    .D(_00428_),
    .Q(\cur_mb_mem[34][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19131_ (.CLK(clknet_leaf_151_clk),
    .D(_00429_),
    .Q(\cur_mb_mem[34][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19132_ (.CLK(clknet_leaf_48_clk),
    .D(_00430_),
    .Q(\cur_mb_mem[34][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19133_ (.CLK(clknet_leaf_247_clk),
    .D(_00431_),
    .Q(\cur_mb_mem[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19134_ (.CLK(clknet_leaf_248_clk),
    .D(_00432_),
    .Q(\cur_mb_mem[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19135_ (.CLK(clknet_leaf_236_clk),
    .D(_00433_),
    .Q(\cur_mb_mem[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19136_ (.CLK(clknet_leaf_248_clk),
    .D(_00434_),
    .Q(\cur_mb_mem[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19137_ (.CLK(clknet_leaf_44_clk),
    .D(_00435_),
    .Q(\cur_mb_mem[35][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19138_ (.CLK(clknet_leaf_58_clk),
    .D(_00436_),
    .Q(\cur_mb_mem[35][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19139_ (.CLK(clknet_leaf_154_clk),
    .D(_00437_),
    .Q(\cur_mb_mem[35][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19140_ (.CLK(clknet_leaf_155_clk),
    .D(_00438_),
    .Q(\cur_mb_mem[35][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19141_ (.CLK(clknet_leaf_65_clk),
    .D(_00439_),
    .Q(\cur_mb_mem[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19142_ (.CLK(clknet_leaf_233_clk),
    .D(_00440_),
    .Q(\cur_mb_mem[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19143_ (.CLK(clknet_leaf_142_clk),
    .D(_00441_),
    .Q(\cur_mb_mem[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19144_ (.CLK(clknet_leaf_64_clk),
    .D(_00442_),
    .Q(\cur_mb_mem[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19145_ (.CLK(clknet_leaf_196_clk),
    .D(_00443_),
    .Q(\cur_mb_mem[36][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19146_ (.CLK(clknet_leaf_195_clk),
    .D(_00444_),
    .Q(\cur_mb_mem[36][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19147_ (.CLK(clknet_leaf_42_clk),
    .D(_00445_),
    .Q(\cur_mb_mem[36][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19148_ (.CLK(clknet_leaf_240_clk),
    .D(_00446_),
    .Q(\cur_mb_mem[36][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19149_ (.CLK(clknet_leaf_257_clk),
    .D(_00447_),
    .Q(\cur_mb_mem[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19150_ (.CLK(clknet_leaf_254_clk),
    .D(_00448_),
    .Q(\cur_mb_mem[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19151_ (.CLK(clknet_leaf_257_clk),
    .D(_00449_),
    .Q(\cur_mb_mem[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19152_ (.CLK(clknet_leaf_257_clk),
    .D(_00450_),
    .Q(\cur_mb_mem[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19153_ (.CLK(clknet_leaf_252_clk),
    .D(_00451_),
    .Q(\cur_mb_mem[37][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19154_ (.CLK(clknet_leaf_252_clk),
    .D(_00452_),
    .Q(\cur_mb_mem[37][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19155_ (.CLK(clknet_leaf_319_clk),
    .D(_00453_),
    .Q(\cur_mb_mem[37][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19156_ (.CLK(clknet_leaf_251_clk),
    .D(_00454_),
    .Q(\cur_mb_mem[37][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19157_ (.CLK(clknet_leaf_227_clk),
    .D(_00455_),
    .Q(\cur_mb_mem[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19158_ (.CLK(clknet_leaf_249_clk),
    .D(_00456_),
    .Q(\cur_mb_mem[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19159_ (.CLK(clknet_leaf_227_clk),
    .D(_00457_),
    .Q(\cur_mb_mem[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19160_ (.CLK(clknet_leaf_227_clk),
    .D(_00458_),
    .Q(\cur_mb_mem[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19161_ (.CLK(clknet_leaf_261_clk),
    .D(_00459_),
    .Q(\cur_mb_mem[38][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19162_ (.CLK(clknet_leaf_262_clk),
    .D(_00460_),
    .Q(\cur_mb_mem[38][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19163_ (.CLK(clknet_leaf_244_clk),
    .D(_00461_),
    .Q(\cur_mb_mem[38][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19164_ (.CLK(clknet_leaf_245_clk),
    .D(_00462_),
    .Q(\cur_mb_mem[38][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19165_ (.CLK(clknet_leaf_261_clk),
    .D(_00463_),
    .Q(\cur_mb_mem[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19166_ (.CLK(clknet_leaf_250_clk),
    .D(_00464_),
    .Q(\cur_mb_mem[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19167_ (.CLK(clknet_leaf_260_clk),
    .D(_00465_),
    .Q(\cur_mb_mem[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19168_ (.CLK(clknet_leaf_261_clk),
    .D(_00466_),
    .Q(\cur_mb_mem[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19169_ (.CLK(clknet_leaf_249_clk),
    .D(_00467_),
    .Q(\cur_mb_mem[39][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19170_ (.CLK(clknet_leaf_261_clk),
    .D(_00468_),
    .Q(\cur_mb_mem[39][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19171_ (.CLK(clknet_leaf_251_clk),
    .D(_00469_),
    .Q(\cur_mb_mem[39][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19172_ (.CLK(clknet_leaf_245_clk),
    .D(_00470_),
    .Q(\cur_mb_mem[39][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19173_ (.CLK(clknet_leaf_33_clk),
    .D(_00471_),
    .Q(\cur_mb_mem[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19174_ (.CLK(clknet_leaf_54_clk),
    .D(_00472_),
    .Q(\cur_mb_mem[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19175_ (.CLK(clknet_leaf_33_clk),
    .D(_00473_),
    .Q(\cur_mb_mem[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19176_ (.CLK(clknet_leaf_29_clk),
    .D(_00474_),
    .Q(\cur_mb_mem[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19177_ (.CLK(clknet_leaf_108_clk),
    .D(_00475_),
    .Q(\cur_mb_mem[40][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19178_ (.CLK(clknet_leaf_108_clk),
    .D(_00476_),
    .Q(\cur_mb_mem[40][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19179_ (.CLK(clknet_leaf_329_clk),
    .D(_00477_),
    .Q(\cur_mb_mem[40][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19180_ (.CLK(clknet_leaf_47_clk),
    .D(_00478_),
    .Q(\cur_mb_mem[40][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19181_ (.CLK(clknet_leaf_253_clk),
    .D(_00479_),
    .Q(\cur_mb_mem[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19182_ (.CLK(clknet_leaf_32_clk),
    .D(_00480_),
    .Q(\cur_mb_mem[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19183_ (.CLK(clknet_leaf_234_clk),
    .D(_00481_),
    .Q(\cur_mb_mem[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19184_ (.CLK(clknet_leaf_249_clk),
    .D(_00482_),
    .Q(\cur_mb_mem[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19185_ (.CLK(clknet_leaf_14_clk),
    .D(_00483_),
    .Q(\cur_mb_mem[41][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19186_ (.CLK(clknet_leaf_14_clk),
    .D(_00484_),
    .Q(\cur_mb_mem[41][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19187_ (.CLK(clknet_leaf_153_clk),
    .D(_00485_),
    .Q(\cur_mb_mem[41][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19188_ (.CLK(clknet_leaf_340_clk),
    .D(_00486_),
    .Q(\cur_mb_mem[41][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19189_ (.CLK(clknet_leaf_70_clk),
    .D(_00487_),
    .Q(\cur_mb_mem[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19190_ (.CLK(clknet_leaf_40_clk),
    .D(_00488_),
    .Q(\cur_mb_mem[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19191_ (.CLK(clknet_leaf_69_clk),
    .D(_00489_),
    .Q(\cur_mb_mem[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19192_ (.CLK(clknet_leaf_66_clk),
    .D(_00490_),
    .Q(\cur_mb_mem[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19193_ (.CLK(clknet_leaf_11_clk),
    .D(_00491_),
    .Q(\cur_mb_mem[42][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19194_ (.CLK(clknet_leaf_12_clk),
    .D(_00492_),
    .Q(\cur_mb_mem[42][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19195_ (.CLK(clknet_leaf_18_clk),
    .D(_00493_),
    .Q(\cur_mb_mem[42][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19196_ (.CLK(clknet_leaf_40_clk),
    .D(_00494_),
    .Q(\cur_mb_mem[42][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19197_ (.CLK(clknet_leaf_67_clk),
    .D(_00495_),
    .Q(\cur_mb_mem[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19198_ (.CLK(clknet_leaf_36_clk),
    .D(_00496_),
    .Q(\cur_mb_mem[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19199_ (.CLK(clknet_leaf_94_clk),
    .D(_00497_),
    .Q(\cur_mb_mem[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19200_ (.CLK(clknet_leaf_65_clk),
    .D(_00498_),
    .Q(\cur_mb_mem[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19201_ (.CLK(clknet_leaf_16_clk),
    .D(_00499_),
    .Q(\cur_mb_mem[43][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19202_ (.CLK(clknet_leaf_18_clk),
    .D(_00500_),
    .Q(\cur_mb_mem[43][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19203_ (.CLK(clknet_leaf_39_clk),
    .D(_00501_),
    .Q(\cur_mb_mem[43][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19204_ (.CLK(clknet_leaf_138_clk),
    .D(_00502_),
    .Q(\cur_mb_mem[43][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19205_ (.CLK(clknet_leaf_141_clk),
    .D(_00503_),
    .Q(\cur_mb_mem[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19206_ (.CLK(clknet_leaf_232_clk),
    .D(_00504_),
    .Q(\cur_mb_mem[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19207_ (.CLK(clknet_leaf_139_clk),
    .D(_00505_),
    .Q(\cur_mb_mem[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19208_ (.CLK(clknet_leaf_140_clk),
    .D(_00506_),
    .Q(\cur_mb_mem[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19209_ (.CLK(clknet_leaf_191_clk),
    .D(_00507_),
    .Q(\cur_mb_mem[44][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19210_ (.CLK(clknet_leaf_192_clk),
    .D(_00508_),
    .Q(\cur_mb_mem[44][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19211_ (.CLK(clknet_leaf_333_clk),
    .D(_00509_),
    .Q(\cur_mb_mem[44][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19212_ (.CLK(clknet_leaf_47_clk),
    .D(_00510_),
    .Q(\cur_mb_mem[44][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19213_ (.CLK(clknet_leaf_169_clk),
    .D(_00511_),
    .Q(\cur_mb_mem[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19214_ (.CLK(clknet_leaf_163_clk),
    .D(_00512_),
    .Q(\cur_mb_mem[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19215_ (.CLK(clknet_leaf_167_clk),
    .D(_00513_),
    .Q(\cur_mb_mem[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19216_ (.CLK(clknet_leaf_169_clk),
    .D(_00514_),
    .Q(\cur_mb_mem[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19217_ (.CLK(clknet_leaf_103_clk),
    .D(_00515_),
    .Q(\cur_mb_mem[45][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19218_ (.CLK(clknet_leaf_104_clk),
    .D(_00516_),
    .Q(\cur_mb_mem[45][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19219_ (.CLK(clknet_leaf_158_clk),
    .D(_00517_),
    .Q(\cur_mb_mem[45][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19220_ (.CLK(clknet_leaf_142_clk),
    .D(_00518_),
    .Q(\cur_mb_mem[45][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19221_ (.CLK(clknet_leaf_195_clk),
    .D(_00519_),
    .Q(\cur_mb_mem[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19222_ (.CLK(clknet_leaf_236_clk),
    .D(_00520_),
    .Q(\cur_mb_mem[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19223_ (.CLK(clknet_leaf_168_clk),
    .D(_00521_),
    .Q(\cur_mb_mem[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19224_ (.CLK(clknet_leaf_193_clk),
    .D(_00522_),
    .Q(\cur_mb_mem[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19225_ (.CLK(clknet_leaf_103_clk),
    .D(_00523_),
    .Q(\cur_mb_mem[46][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19226_ (.CLK(clknet_leaf_107_clk),
    .D(_00524_),
    .Q(\cur_mb_mem[46][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19227_ (.CLK(clknet_leaf_328_clk),
    .D(_00525_),
    .Q(\cur_mb_mem[46][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19228_ (.CLK(clknet_leaf_328_clk),
    .D(_00526_),
    .Q(\cur_mb_mem[46][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19229_ (.CLK(clknet_leaf_93_clk),
    .D(_00527_),
    .Q(\cur_mb_mem[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19230_ (.CLK(clknet_leaf_233_clk),
    .D(_00528_),
    .Q(\cur_mb_mem[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19231_ (.CLK(clknet_leaf_63_clk),
    .D(_00529_),
    .Q(\cur_mb_mem[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19232_ (.CLK(clknet_leaf_93_clk),
    .D(_00530_),
    .Q(\cur_mb_mem[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19233_ (.CLK(clknet_leaf_134_clk),
    .D(_00531_),
    .Q(\cur_mb_mem[47][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19234_ (.CLK(clknet_leaf_134_clk),
    .D(_00532_),
    .Q(\cur_mb_mem[47][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19235_ (.CLK(clknet_leaf_244_clk),
    .D(_00533_),
    .Q(\cur_mb_mem[47][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19236_ (.CLK(clknet_leaf_251_clk),
    .D(_00534_),
    .Q(\cur_mb_mem[47][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19237_ (.CLK(clknet_leaf_250_clk),
    .D(_00535_),
    .Q(\cur_mb_mem[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19238_ (.CLK(clknet_leaf_172_clk),
    .D(_00536_),
    .Q(\cur_mb_mem[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19239_ (.CLK(clknet_leaf_234_clk),
    .D(_00537_),
    .Q(\cur_mb_mem[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19240_ (.CLK(clknet_leaf_250_clk),
    .D(_00538_),
    .Q(\cur_mb_mem[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19241_ (.CLK(clknet_leaf_113_clk),
    .D(_00539_),
    .Q(\cur_mb_mem[48][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19242_ (.CLK(clknet_leaf_113_clk),
    .D(_00540_),
    .Q(\cur_mb_mem[48][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19243_ (.CLK(clknet_leaf_165_clk),
    .D(_00541_),
    .Q(\cur_mb_mem[48][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19244_ (.CLK(clknet_leaf_144_clk),
    .D(_00542_),
    .Q(\cur_mb_mem[48][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19245_ (.CLK(clknet_leaf_247_clk),
    .D(_00543_),
    .Q(\cur_mb_mem[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19246_ (.CLK(clknet_leaf_171_clk),
    .D(_00544_),
    .Q(\cur_mb_mem[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19247_ (.CLK(clknet_leaf_234_clk),
    .D(_00545_),
    .Q(\cur_mb_mem[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19248_ (.CLK(clknet_leaf_235_clk),
    .D(_00546_),
    .Q(\cur_mb_mem[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19249_ (.CLK(clknet_leaf_195_clk),
    .D(_00547_),
    .Q(\cur_mb_mem[49][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19250_ (.CLK(clknet_leaf_194_clk),
    .D(_00548_),
    .Q(\cur_mb_mem[49][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19251_ (.CLK(clknet_leaf_162_clk),
    .D(_00549_),
    .Q(\cur_mb_mem[49][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19252_ (.CLK(clknet_leaf_236_clk),
    .D(_00550_),
    .Q(\cur_mb_mem[49][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19253_ (.CLK(clknet_leaf_316_clk),
    .D(_00551_),
    .Q(\cur_mb_mem[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19254_ (.CLK(clknet_leaf_193_clk),
    .D(_00552_),
    .Q(\cur_mb_mem[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19255_ (.CLK(clknet_leaf_316_clk),
    .D(_00553_),
    .Q(\cur_mb_mem[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19256_ (.CLK(clknet_leaf_317_clk),
    .D(_00554_),
    .Q(\cur_mb_mem[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19257_ (.CLK(clknet_leaf_194_clk),
    .D(_00555_),
    .Q(\cur_mb_mem[50][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19258_ (.CLK(clknet_leaf_195_clk),
    .D(_00556_),
    .Q(\cur_mb_mem[50][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19259_ (.CLK(clknet_leaf_170_clk),
    .D(_00557_),
    .Q(\cur_mb_mem[50][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19260_ (.CLK(clknet_leaf_245_clk),
    .D(_00558_),
    .Q(\cur_mb_mem[50][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19261_ (.CLK(clknet_leaf_227_clk),
    .D(_00559_),
    .Q(\cur_mb_mem[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19262_ (.CLK(clknet_leaf_224_clk),
    .D(_00560_),
    .Q(\cur_mb_mem[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19263_ (.CLK(clknet_leaf_162_clk),
    .D(_00561_),
    .Q(\cur_mb_mem[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19264_ (.CLK(clknet_leaf_228_clk),
    .D(_00562_),
    .Q(\cur_mb_mem[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19265_ (.CLK(clknet_leaf_263_clk),
    .D(_00563_),
    .Q(\cur_mb_mem[51][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19266_ (.CLK(clknet_leaf_224_clk),
    .D(_00564_),
    .Q(\cur_mb_mem[51][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19267_ (.CLK(clknet_leaf_239_clk),
    .D(_00565_),
    .Q(\cur_mb_mem[51][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19268_ (.CLK(clknet_leaf_239_clk),
    .D(_00566_),
    .Q(\cur_mb_mem[51][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19269_ (.CLK(clknet_leaf_89_clk),
    .D(_00567_),
    .Q(\cur_mb_mem[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19270_ (.CLK(clknet_leaf_127_clk),
    .D(_00568_),
    .Q(\cur_mb_mem[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19271_ (.CLK(clknet_leaf_89_clk),
    .D(_00569_),
    .Q(\cur_mb_mem[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19272_ (.CLK(clknet_leaf_91_clk),
    .D(_00570_),
    .Q(\cur_mb_mem[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19273_ (.CLK(clknet_leaf_194_clk),
    .D(_00571_),
    .Q(\cur_mb_mem[52][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19274_ (.CLK(clknet_leaf_194_clk),
    .D(_00572_),
    .Q(\cur_mb_mem[52][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19275_ (.CLK(clknet_leaf_158_clk),
    .D(_00573_),
    .Q(\cur_mb_mem[52][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19276_ (.CLK(clknet_leaf_147_clk),
    .D(_00574_),
    .Q(\cur_mb_mem[52][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19277_ (.CLK(clknet_leaf_273_clk),
    .D(_00575_),
    .Q(\cur_mb_mem[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19278_ (.CLK(clknet_leaf_321_clk),
    .D(_00576_),
    .Q(\cur_mb_mem[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19279_ (.CLK(clknet_leaf_315_clk),
    .D(_00577_),
    .Q(\cur_mb_mem[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19280_ (.CLK(clknet_leaf_282_clk),
    .D(_00578_),
    .Q(\cur_mb_mem[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19281_ (.CLK(clknet_leaf_228_clk),
    .D(_00579_),
    .Q(\cur_mb_mem[53][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19282_ (.CLK(clknet_leaf_196_clk),
    .D(_00580_),
    .Q(\cur_mb_mem[53][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19283_ (.CLK(clknet_leaf_175_clk),
    .D(_00581_),
    .Q(\cur_mb_mem[53][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19284_ (.CLK(clknet_leaf_307_clk),
    .D(_00582_),
    .Q(\cur_mb_mem[53][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19285_ (.CLK(clknet_leaf_262_clk),
    .D(_00583_),
    .Q(\cur_mb_mem[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19286_ (.CLK(clknet_leaf_224_clk),
    .D(_00584_),
    .Q(\cur_mb_mem[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19287_ (.CLK(clknet_leaf_234_clk),
    .D(_00585_),
    .Q(\cur_mb_mem[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19288_ (.CLK(clknet_leaf_263_clk),
    .D(_00586_),
    .Q(\cur_mb_mem[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19289_ (.CLK(clknet_leaf_220_clk),
    .D(_00587_),
    .Q(\cur_mb_mem[54][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19290_ (.CLK(clknet_leaf_220_clk),
    .D(_00588_),
    .Q(\cur_mb_mem[54][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19291_ (.CLK(clknet_leaf_162_clk),
    .D(_00589_),
    .Q(\cur_mb_mem[54][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19292_ (.CLK(clknet_leaf_327_clk),
    .D(_00590_),
    .Q(\cur_mb_mem[54][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19293_ (.CLK(clknet_leaf_257_clk),
    .D(_00591_),
    .Q(\cur_mb_mem[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19294_ (.CLK(clknet_leaf_254_clk),
    .D(_00592_),
    .Q(\cur_mb_mem[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19295_ (.CLK(clknet_leaf_250_clk),
    .D(_00593_),
    .Q(\cur_mb_mem[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19296_ (.CLK(clknet_leaf_260_clk),
    .D(_00594_),
    .Q(\cur_mb_mem[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19297_ (.CLK(clknet_leaf_226_clk),
    .D(_00595_),
    .Q(\cur_mb_mem[55][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19298_ (.CLK(clknet_leaf_226_clk),
    .D(_00596_),
    .Q(\cur_mb_mem[55][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19299_ (.CLK(clknet_leaf_313_clk),
    .D(_00597_),
    .Q(\cur_mb_mem[55][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19300_ (.CLK(clknet_leaf_251_clk),
    .D(_00598_),
    .Q(\cur_mb_mem[55][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19301_ (.CLK(clknet_leaf_315_clk),
    .D(_00599_),
    .Q(\cur_mb_mem[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19302_ (.CLK(clknet_leaf_232_clk),
    .D(_00600_),
    .Q(\cur_mb_mem[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19303_ (.CLK(clknet_leaf_315_clk),
    .D(_00601_),
    .Q(\cur_mb_mem[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19304_ (.CLK(clknet_leaf_254_clk),
    .D(_00602_),
    .Q(\cur_mb_mem[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19305_ (.CLK(clknet_leaf_192_clk),
    .D(_00603_),
    .Q(\cur_mb_mem[56][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19306_ (.CLK(clknet_leaf_193_clk),
    .D(_00604_),
    .Q(\cur_mb_mem[56][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19307_ (.CLK(clknet_leaf_232_clk),
    .D(_00605_),
    .Q(\cur_mb_mem[56][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19308_ (.CLK(clknet_leaf_245_clk),
    .D(_00606_),
    .Q(\cur_mb_mem[56][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19309_ (.CLK(clknet_leaf_112_clk),
    .D(_00607_),
    .Q(\cur_mb_mem[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19310_ (.CLK(clknet_leaf_127_clk),
    .D(_00608_),
    .Q(\cur_mb_mem[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19311_ (.CLK(clknet_leaf_131_clk),
    .D(_00609_),
    .Q(\cur_mb_mem[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19312_ (.CLK(clknet_leaf_112_clk),
    .D(_00610_),
    .Q(\cur_mb_mem[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19313_ (.CLK(clknet_leaf_171_clk),
    .D(_00611_),
    .Q(\cur_mb_mem[57][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19314_ (.CLK(clknet_leaf_168_clk),
    .D(_00612_),
    .Q(\cur_mb_mem[57][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19315_ (.CLK(clknet_leaf_239_clk),
    .D(_00613_),
    .Q(\cur_mb_mem[57][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19316_ (.CLK(clknet_leaf_150_clk),
    .D(_00614_),
    .Q(\cur_mb_mem[57][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19317_ (.CLK(clknet_leaf_179_clk),
    .D(_00615_),
    .Q(\cur_mb_mem[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19318_ (.CLK(clknet_leaf_325_clk),
    .D(_00616_),
    .Q(\cur_mb_mem[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19319_ (.CLK(clknet_leaf_142_clk),
    .D(_00617_),
    .Q(\cur_mb_mem[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19320_ (.CLK(clknet_leaf_134_clk),
    .D(_00618_),
    .Q(\cur_mb_mem[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19321_ (.CLK(clknet_leaf_133_clk),
    .D(_00619_),
    .Q(\cur_mb_mem[58][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19322_ (.CLK(clknet_leaf_132_clk),
    .D(_00620_),
    .Q(\cur_mb_mem[58][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19323_ (.CLK(clknet_leaf_337_clk),
    .D(_00621_),
    .Q(\cur_mb_mem[58][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19324_ (.CLK(clknet_leaf_53_clk),
    .D(_00622_),
    .Q(\cur_mb_mem[58][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19325_ (.CLK(clknet_leaf_317_clk),
    .D(_00623_),
    .Q(\cur_mb_mem[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19326_ (.CLK(clknet_leaf_326_clk),
    .D(_00624_),
    .Q(\cur_mb_mem[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19327_ (.CLK(clknet_leaf_317_clk),
    .D(_00625_),
    .Q(\cur_mb_mem[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19328_ (.CLK(clknet_leaf_318_clk),
    .D(_00626_),
    .Q(\cur_mb_mem[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19329_ (.CLK(clknet_leaf_255_clk),
    .D(_00627_),
    .Q(\cur_mb_mem[59][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19330_ (.CLK(clknet_leaf_256_clk),
    .D(_00628_),
    .Q(\cur_mb_mem[59][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19331_ (.CLK(clknet_leaf_327_clk),
    .D(_00629_),
    .Q(\cur_mb_mem[59][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19332_ (.CLK(clknet_leaf_239_clk),
    .D(_00630_),
    .Q(\cur_mb_mem[59][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19333_ (.CLK(clknet_leaf_273_clk),
    .D(_00631_),
    .Q(\cur_mb_mem[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19334_ (.CLK(clknet_leaf_243_clk),
    .D(_00632_),
    .Q(\cur_mb_mem[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19335_ (.CLK(clknet_leaf_315_clk),
    .D(_00633_),
    .Q(\cur_mb_mem[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19336_ (.CLK(clknet_leaf_248_clk),
    .D(_00634_),
    .Q(\cur_mb_mem[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19337_ (.CLK(clknet_leaf_226_clk),
    .D(_00635_),
    .Q(\cur_mb_mem[60][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19338_ (.CLK(clknet_leaf_226_clk),
    .D(_00636_),
    .Q(\cur_mb_mem[60][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19339_ (.CLK(clknet_leaf_53_clk),
    .D(_00637_),
    .Q(\cur_mb_mem[60][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19340_ (.CLK(clknet_leaf_342_clk),
    .D(_00638_),
    .Q(\cur_mb_mem[60][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19341_ (.CLK(clknet_leaf_95_clk),
    .D(_00639_),
    .Q(\cur_mb_mem[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19342_ (.CLK(clknet_leaf_236_clk),
    .D(_00640_),
    .Q(\cur_mb_mem[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19343_ (.CLK(clknet_leaf_94_clk),
    .D(_00641_),
    .Q(\cur_mb_mem[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19344_ (.CLK(clknet_leaf_65_clk),
    .D(_00642_),
    .Q(\cur_mb_mem[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19345_ (.CLK(clknet_leaf_192_clk),
    .D(_00643_),
    .Q(\cur_mb_mem[61][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19346_ (.CLK(clknet_leaf_192_clk),
    .D(_00644_),
    .Q(\cur_mb_mem[61][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19347_ (.CLK(clknet_leaf_72_clk),
    .D(_00645_),
    .Q(\cur_mb_mem[61][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19348_ (.CLK(clknet_leaf_240_clk),
    .D(_00646_),
    .Q(\cur_mb_mem[61][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19349_ (.CLK(clknet_leaf_179_clk),
    .D(_00647_),
    .Q(\cur_mb_mem[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19350_ (.CLK(clknet_leaf_172_clk),
    .D(_00648_),
    .Q(\cur_mb_mem[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19351_ (.CLK(clknet_leaf_174_clk),
    .D(_00649_),
    .Q(\cur_mb_mem[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19352_ (.CLK(clknet_leaf_127_clk),
    .D(_00650_),
    .Q(\cur_mb_mem[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19353_ (.CLK(clknet_leaf_133_clk),
    .D(_00651_),
    .Q(\cur_mb_mem[62][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19354_ (.CLK(clknet_leaf_133_clk),
    .D(_00652_),
    .Q(\cur_mb_mem[62][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19355_ (.CLK(clknet_leaf_337_clk),
    .D(_00653_),
    .Q(\cur_mb_mem[62][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19356_ (.CLK(clknet_leaf_242_clk),
    .D(_00654_),
    .Q(\cur_mb_mem[62][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19357_ (.CLK(clknet_leaf_254_clk),
    .D(_00655_),
    .Q(\cur_mb_mem[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19358_ (.CLK(clknet_leaf_317_clk),
    .D(_00656_),
    .Q(\cur_mb_mem[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19359_ (.CLK(clknet_leaf_255_clk),
    .D(_00657_),
    .Q(\cur_mb_mem[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19360_ (.CLK(clknet_leaf_250_clk),
    .D(_00658_),
    .Q(\cur_mb_mem[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19361_ (.CLK(clknet_leaf_255_clk),
    .D(_00659_),
    .Q(\cur_mb_mem[63][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19362_ (.CLK(clknet_leaf_255_clk),
    .D(_00660_),
    .Q(\cur_mb_mem[63][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19363_ (.CLK(clknet_leaf_318_clk),
    .D(_00661_),
    .Q(\cur_mb_mem[63][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19364_ (.CLK(clknet_leaf_245_clk),
    .D(_00662_),
    .Q(\cur_mb_mem[63][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19365_ (.CLK(clknet_leaf_136_clk),
    .D(_00663_),
    .Q(\cur_mb_mem[64][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19366_ (.CLK(clknet_leaf_129_clk),
    .D(_00664_),
    .Q(\cur_mb_mem[64][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19367_ (.CLK(clknet_leaf_131_clk),
    .D(_00665_),
    .Q(\cur_mb_mem[64][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19368_ (.CLK(clknet_leaf_115_clk),
    .D(_00666_),
    .Q(\cur_mb_mem[64][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19369_ (.CLK(clknet_leaf_114_clk),
    .D(_00667_),
    .Q(\cur_mb_mem[64][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19370_ (.CLK(clknet_leaf_113_clk),
    .D(_00668_),
    .Q(\cur_mb_mem[64][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19371_ (.CLK(clknet_leaf_161_clk),
    .D(_00669_),
    .Q(\cur_mb_mem[64][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19372_ (.CLK(clknet_leaf_162_clk),
    .D(_00670_),
    .Q(\cur_mb_mem[64][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19373_ (.CLK(clknet_leaf_108_clk),
    .D(_00671_),
    .Q(\cur_mb_mem[65][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19374_ (.CLK(clknet_leaf_137_clk),
    .D(_00672_),
    .Q(\cur_mb_mem[65][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19375_ (.CLK(clknet_leaf_112_clk),
    .D(_00673_),
    .Q(\cur_mb_mem[65][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19376_ (.CLK(clknet_leaf_115_clk),
    .D(_00674_),
    .Q(\cur_mb_mem[65][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19377_ (.CLK(clknet_leaf_114_clk),
    .D(_00675_),
    .Q(\cur_mb_mem[65][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19378_ (.CLK(clknet_leaf_119_clk),
    .D(_00676_),
    .Q(\cur_mb_mem[65][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19379_ (.CLK(clknet_leaf_138_clk),
    .D(_00677_),
    .Q(\cur_mb_mem[65][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19380_ (.CLK(clknet_leaf_139_clk),
    .D(_00678_),
    .Q(\cur_mb_mem[65][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19381_ (.CLK(clknet_leaf_88_clk),
    .D(_00679_),
    .Q(\cur_mb_mem[66][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19382_ (.CLK(clknet_leaf_137_clk),
    .D(_00680_),
    .Q(\cur_mb_mem[66][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19383_ (.CLK(clknet_leaf_101_clk),
    .D(_00681_),
    .Q(\cur_mb_mem[66][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19384_ (.CLK(clknet_leaf_99_clk),
    .D(_00682_),
    .Q(\cur_mb_mem[66][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19385_ (.CLK(clknet_leaf_117_clk),
    .D(_00683_),
    .Q(\cur_mb_mem[66][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19386_ (.CLK(clknet_leaf_117_clk),
    .D(_00684_),
    .Q(\cur_mb_mem[66][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19387_ (.CLK(clknet_leaf_176_clk),
    .D(_00685_),
    .Q(\cur_mb_mem[66][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19388_ (.CLK(clknet_leaf_176_clk),
    .D(_00686_),
    .Q(\cur_mb_mem[66][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19389_ (.CLK(clknet_leaf_101_clk),
    .D(_00687_),
    .Q(\cur_mb_mem[67][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19390_ (.CLK(clknet_leaf_137_clk),
    .D(_00688_),
    .Q(\cur_mb_mem[67][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19391_ (.CLK(clknet_leaf_100_clk),
    .D(_00689_),
    .Q(\cur_mb_mem[67][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19392_ (.CLK(clknet_leaf_98_clk),
    .D(_00690_),
    .Q(\cur_mb_mem[67][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19393_ (.CLK(clknet_leaf_117_clk),
    .D(_00691_),
    .Q(\cur_mb_mem[67][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19394_ (.CLK(clknet_leaf_117_clk),
    .D(_00692_),
    .Q(\cur_mb_mem[67][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19395_ (.CLK(clknet_leaf_130_clk),
    .D(_00693_),
    .Q(\cur_mb_mem[67][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19396_ (.CLK(clknet_leaf_131_clk),
    .D(_00694_),
    .Q(\cur_mb_mem[67][7] ));
 sky130_fd_sc_hd__dfxtp_2 _19397_ (.CLK(clknet_leaf_95_clk),
    .D(_00695_),
    .Q(\cur_mb_mem[68][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19398_ (.CLK(clknet_leaf_138_clk),
    .D(_00696_),
    .Q(\cur_mb_mem[68][1] ));
 sky130_fd_sc_hd__dfxtp_2 _19399_ (.CLK(clknet_leaf_95_clk),
    .D(_00697_),
    .Q(\cur_mb_mem[68][2] ));
 sky130_fd_sc_hd__dfxtp_4 _19400_ (.CLK(clknet_leaf_103_clk),
    .D(_00698_),
    .Q(\cur_mb_mem[68][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19401_ (.CLK(clknet_leaf_102_clk),
    .D(_00699_),
    .Q(\cur_mb_mem[68][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19402_ (.CLK(clknet_leaf_102_clk),
    .D(_00700_),
    .Q(\cur_mb_mem[68][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19403_ (.CLK(clknet_leaf_138_clk),
    .D(_00701_),
    .Q(\cur_mb_mem[68][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19404_ (.CLK(clknet_leaf_139_clk),
    .D(_00702_),
    .Q(\cur_mb_mem[68][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19405_ (.CLK(clknet_leaf_108_clk),
    .D(_00703_),
    .Q(\cur_mb_mem[69][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19406_ (.CLK(clknet_leaf_130_clk),
    .D(_00704_),
    .Q(\cur_mb_mem[69][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19407_ (.CLK(clknet_leaf_135_clk),
    .D(_00705_),
    .Q(\cur_mb_mem[69][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19408_ (.CLK(clknet_leaf_115_clk),
    .D(_00706_),
    .Q(\cur_mb_mem[69][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19409_ (.CLK(clknet_leaf_102_clk),
    .D(_00707_),
    .Q(\cur_mb_mem[69][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19410_ (.CLK(clknet_leaf_102_clk),
    .D(_00708_),
    .Q(\cur_mb_mem[69][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19411_ (.CLK(clknet_leaf_130_clk),
    .D(_00709_),
    .Q(\cur_mb_mem[69][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19412_ (.CLK(clknet_leaf_130_clk),
    .D(_00710_),
    .Q(\cur_mb_mem[69][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19413_ (.CLK(clknet_leaf_108_clk),
    .D(_00711_),
    .Q(\cur_mb_mem[70][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19414_ (.CLK(clknet_leaf_95_clk),
    .D(_00712_),
    .Q(\cur_mb_mem[70][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19415_ (.CLK(clknet_leaf_112_clk),
    .D(_00713_),
    .Q(\cur_mb_mem[70][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19416_ (.CLK(clknet_leaf_115_clk),
    .D(_00714_),
    .Q(\cur_mb_mem[70][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19417_ (.CLK(clknet_leaf_102_clk),
    .D(_00715_),
    .Q(\cur_mb_mem[70][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19418_ (.CLK(clknet_leaf_102_clk),
    .D(_00716_),
    .Q(\cur_mb_mem[70][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19419_ (.CLK(clknet_leaf_130_clk),
    .D(_00717_),
    .Q(\cur_mb_mem[70][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19420_ (.CLK(clknet_leaf_136_clk),
    .D(_00718_),
    .Q(\cur_mb_mem[70][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19421_ (.CLK(clknet_leaf_97_clk),
    .D(_00719_),
    .Q(\cur_mb_mem[71][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19422_ (.CLK(clknet_leaf_161_clk),
    .D(_00720_),
    .Q(\cur_mb_mem[71][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19423_ (.CLK(clknet_leaf_64_clk),
    .D(_00721_),
    .Q(\cur_mb_mem[71][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19424_ (.CLK(clknet_leaf_105_clk),
    .D(_00722_),
    .Q(\cur_mb_mem[71][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19425_ (.CLK(clknet_leaf_114_clk),
    .D(_00723_),
    .Q(\cur_mb_mem[71][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19426_ (.CLK(clknet_leaf_113_clk),
    .D(_00724_),
    .Q(\cur_mb_mem[71][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19427_ (.CLK(clknet_leaf_160_clk),
    .D(_00725_),
    .Q(\cur_mb_mem[71][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19428_ (.CLK(clknet_leaf_161_clk),
    .D(_00726_),
    .Q(\cur_mb_mem[71][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19429_ (.CLK(clknet_leaf_88_clk),
    .D(_00727_),
    .Q(\cur_mb_mem[72][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19430_ (.CLK(clknet_leaf_135_clk),
    .D(_00728_),
    .Q(\cur_mb_mem[72][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19431_ (.CLK(clknet_leaf_88_clk),
    .D(_00729_),
    .Q(\cur_mb_mem[72][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19432_ (.CLK(clknet_leaf_105_clk),
    .D(_00730_),
    .Q(\cur_mb_mem[72][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19433_ (.CLK(clknet_leaf_118_clk),
    .D(_00731_),
    .Q(\cur_mb_mem[72][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19434_ (.CLK(clknet_leaf_118_clk),
    .D(_00732_),
    .Q(\cur_mb_mem[72][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19435_ (.CLK(clknet_leaf_145_clk),
    .D(_00733_),
    .Q(\cur_mb_mem[72][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19436_ (.CLK(clknet_leaf_129_clk),
    .D(_00734_),
    .Q(\cur_mb_mem[72][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19437_ (.CLK(clknet_leaf_101_clk),
    .D(_00735_),
    .Q(\cur_mb_mem[73][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19438_ (.CLK(clknet_leaf_64_clk),
    .D(_00736_),
    .Q(\cur_mb_mem[73][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19439_ (.CLK(clknet_leaf_101_clk),
    .D(_00737_),
    .Q(\cur_mb_mem[73][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19440_ (.CLK(clknet_leaf_97_clk),
    .D(_00738_),
    .Q(\cur_mb_mem[73][3] ));
 sky130_fd_sc_hd__dfxtp_2 _19441_ (.CLK(clknet_leaf_134_clk),
    .D(_00739_),
    .Q(\cur_mb_mem[73][4] ));
 sky130_fd_sc_hd__dfxtp_2 _19442_ (.CLK(clknet_leaf_136_clk),
    .D(_00740_),
    .Q(\cur_mb_mem[73][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19443_ (.CLK(clknet_leaf_138_clk),
    .D(_00741_),
    .Q(\cur_mb_mem[73][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19444_ (.CLK(clknet_leaf_139_clk),
    .D(_00742_),
    .Q(\cur_mb_mem[73][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19445_ (.CLK(clknet_leaf_96_clk),
    .D(_00743_),
    .Q(\cur_mb_mem[74][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19446_ (.CLK(clknet_leaf_137_clk),
    .D(_00744_),
    .Q(\cur_mb_mem[74][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19447_ (.CLK(clknet_leaf_94_clk),
    .D(_00745_),
    .Q(\cur_mb_mem[74][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19448_ (.CLK(clknet_leaf_96_clk),
    .D(_00746_),
    .Q(\cur_mb_mem[74][3] ));
 sky130_fd_sc_hd__dfxtp_2 _19449_ (.CLK(clknet_leaf_135_clk),
    .D(_00747_),
    .Q(\cur_mb_mem[74][4] ));
 sky130_fd_sc_hd__dfxtp_2 _19450_ (.CLK(clknet_leaf_134_clk),
    .D(_00748_),
    .Q(\cur_mb_mem[74][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19451_ (.CLK(clknet_leaf_159_clk),
    .D(_00749_),
    .Q(\cur_mb_mem[74][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19452_ (.CLK(clknet_leaf_137_clk),
    .D(_00750_),
    .Q(\cur_mb_mem[74][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19453_ (.CLK(clknet_leaf_94_clk),
    .D(_00751_),
    .Q(\cur_mb_mem[75][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19454_ (.CLK(clknet_leaf_144_clk),
    .D(_00752_),
    .Q(\cur_mb_mem[75][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19455_ (.CLK(clknet_leaf_68_clk),
    .D(_00753_),
    .Q(\cur_mb_mem[75][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19456_ (.CLK(clknet_leaf_104_clk),
    .D(_00754_),
    .Q(\cur_mb_mem[75][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19457_ (.CLK(clknet_leaf_124_clk),
    .D(_00755_),
    .Q(\cur_mb_mem[75][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19458_ (.CLK(clknet_leaf_119_clk),
    .D(_00756_),
    .Q(\cur_mb_mem[75][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19459_ (.CLK(clknet_leaf_147_clk),
    .D(_00757_),
    .Q(\cur_mb_mem[75][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19460_ (.CLK(clknet_leaf_60_clk),
    .D(_00758_),
    .Q(\cur_mb_mem[75][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19461_ (.CLK(clknet_leaf_167_clk),
    .D(_00759_),
    .Q(\cur_mb_mem[76][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19462_ (.CLK(clknet_leaf_134_clk),
    .D(_00760_),
    .Q(\cur_mb_mem[76][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19463_ (.CLK(clknet_leaf_231_clk),
    .D(_00761_),
    .Q(\cur_mb_mem[76][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19464_ (.CLK(clknet_leaf_185_clk),
    .D(_00762_),
    .Q(\cur_mb_mem[76][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19465_ (.CLK(clknet_leaf_118_clk),
    .D(_00763_),
    .Q(\cur_mb_mem[76][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19466_ (.CLK(clknet_leaf_114_clk),
    .D(_00764_),
    .Q(\cur_mb_mem[76][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19467_ (.CLK(clknet_leaf_157_clk),
    .D(_00765_),
    .Q(\cur_mb_mem[76][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19468_ (.CLK(clknet_leaf_163_clk),
    .D(_00766_),
    .Q(\cur_mb_mem[76][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19469_ (.CLK(clknet_leaf_112_clk),
    .D(_00767_),
    .Q(\cur_mb_mem[77][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19470_ (.CLK(clknet_leaf_127_clk),
    .D(_00768_),
    .Q(\cur_mb_mem[77][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19471_ (.CLK(clknet_leaf_132_clk),
    .D(_00769_),
    .Q(\cur_mb_mem[77][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19472_ (.CLK(clknet_leaf_114_clk),
    .D(_00770_),
    .Q(\cur_mb_mem[77][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19473_ (.CLK(clknet_leaf_118_clk),
    .D(_00771_),
    .Q(\cur_mb_mem[77][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19474_ (.CLK(clknet_leaf_114_clk),
    .D(_00772_),
    .Q(\cur_mb_mem[77][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19475_ (.CLK(clknet_leaf_144_clk),
    .D(_00773_),
    .Q(\cur_mb_mem[77][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19476_ (.CLK(clknet_leaf_144_clk),
    .D(_00774_),
    .Q(\cur_mb_mem[77][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19477_ (.CLK(clknet_leaf_109_clk),
    .D(_00775_),
    .Q(\cur_mb_mem[78][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19478_ (.CLK(clknet_leaf_124_clk),
    .D(_00776_),
    .Q(\cur_mb_mem[78][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19479_ (.CLK(clknet_leaf_131_clk),
    .D(_00777_),
    .Q(\cur_mb_mem[78][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19480_ (.CLK(clknet_leaf_116_clk),
    .D(_00778_),
    .Q(\cur_mb_mem[78][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19481_ (.CLK(clknet_leaf_124_clk),
    .D(_00779_),
    .Q(\cur_mb_mem[78][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19482_ (.CLK(clknet_leaf_120_clk),
    .D(_00780_),
    .Q(\cur_mb_mem[78][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19483_ (.CLK(clknet_leaf_147_clk),
    .D(_00781_),
    .Q(\cur_mb_mem[78][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19484_ (.CLK(clknet_leaf_148_clk),
    .D(_00782_),
    .Q(\cur_mb_mem[78][7] ));
 sky130_fd_sc_hd__dfxtp_2 _19485_ (.CLK(clknet_leaf_229_clk),
    .D(_00783_),
    .Q(\cur_mb_mem[79][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19486_ (.CLK(clknet_leaf_160_clk),
    .D(_00784_),
    .Q(\cur_mb_mem[79][1] ));
 sky130_fd_sc_hd__dfxtp_2 _19487_ (.CLK(clknet_leaf_167_clk),
    .D(_00785_),
    .Q(\cur_mb_mem[79][2] ));
 sky130_fd_sc_hd__dfxtp_2 _19488_ (.CLK(clknet_leaf_169_clk),
    .D(_00786_),
    .Q(\cur_mb_mem[79][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19489_ (.CLK(clknet_leaf_136_clk),
    .D(_00787_),
    .Q(\cur_mb_mem[79][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19490_ (.CLK(clknet_leaf_110_clk),
    .D(_00788_),
    .Q(\cur_mb_mem[79][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19491_ (.CLK(clknet_leaf_159_clk),
    .D(_00789_),
    .Q(\cur_mb_mem[79][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19492_ (.CLK(clknet_leaf_162_clk),
    .D(_00790_),
    .Q(\cur_mb_mem[79][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19493_ (.CLK(clknet_leaf_179_clk),
    .D(_00791_),
    .Q(\cur_mb_mem[80][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19494_ (.CLK(clknet_leaf_145_clk),
    .D(_00792_),
    .Q(\cur_mb_mem[80][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19495_ (.CLK(clknet_leaf_173_clk),
    .D(_00793_),
    .Q(\cur_mb_mem[80][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19496_ (.CLK(clknet_leaf_124_clk),
    .D(_00794_),
    .Q(\cur_mb_mem[80][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19497_ (.CLK(clknet_leaf_124_clk),
    .D(_00795_),
    .Q(\cur_mb_mem[80][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19498_ (.CLK(clknet_leaf_124_clk),
    .D(_00796_),
    .Q(\cur_mb_mem[80][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19499_ (.CLK(clknet_leaf_142_clk),
    .D(_00797_),
    .Q(\cur_mb_mem[80][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19500_ (.CLK(clknet_leaf_147_clk),
    .D(_00798_),
    .Q(\cur_mb_mem[80][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19501_ (.CLK(clknet_leaf_95_clk),
    .D(_00799_),
    .Q(\cur_mb_mem[81][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19502_ (.CLK(clknet_leaf_127_clk),
    .D(_00800_),
    .Q(\cur_mb_mem[81][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19503_ (.CLK(clknet_leaf_131_clk),
    .D(_00801_),
    .Q(\cur_mb_mem[81][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19504_ (.CLK(clknet_leaf_103_clk),
    .D(_00802_),
    .Q(\cur_mb_mem[81][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19505_ (.CLK(clknet_leaf_104_clk),
    .D(_00803_),
    .Q(\cur_mb_mem[81][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19506_ (.CLK(clknet_leaf_105_clk),
    .D(_00804_),
    .Q(\cur_mb_mem[81][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19507_ (.CLK(clknet_leaf_144_clk),
    .D(_00805_),
    .Q(\cur_mb_mem[81][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19508_ (.CLK(clknet_leaf_60_clk),
    .D(_00806_),
    .Q(\cur_mb_mem[81][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19509_ (.CLK(clknet_leaf_143_clk),
    .D(_00807_),
    .Q(\cur_mb_mem[82][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19510_ (.CLK(clknet_leaf_137_clk),
    .D(_00808_),
    .Q(\cur_mb_mem[82][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19511_ (.CLK(clknet_leaf_139_clk),
    .D(_00809_),
    .Q(\cur_mb_mem[82][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19512_ (.CLK(clknet_leaf_119_clk),
    .D(_00810_),
    .Q(\cur_mb_mem[82][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19513_ (.CLK(clknet_leaf_105_clk),
    .D(_00811_),
    .Q(\cur_mb_mem[82][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19514_ (.CLK(clknet_leaf_105_clk),
    .D(_00812_),
    .Q(\cur_mb_mem[82][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19515_ (.CLK(clknet_leaf_144_clk),
    .D(_00813_),
    .Q(\cur_mb_mem[82][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19516_ (.CLK(clknet_leaf_148_clk),
    .D(_00814_),
    .Q(\cur_mb_mem[82][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19517_ (.CLK(clknet_leaf_100_clk),
    .D(_00815_),
    .Q(\cur_mb_mem[83][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19518_ (.CLK(clknet_leaf_126_clk),
    .D(_00816_),
    .Q(\cur_mb_mem[83][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19519_ (.CLK(clknet_leaf_101_clk),
    .D(_00817_),
    .Q(\cur_mb_mem[83][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19520_ (.CLK(clknet_leaf_97_clk),
    .D(_00818_),
    .Q(\cur_mb_mem[83][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19521_ (.CLK(clknet_leaf_99_clk),
    .D(_00819_),
    .Q(\cur_mb_mem[83][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19522_ (.CLK(clknet_leaf_98_clk),
    .D(_00820_),
    .Q(\cur_mb_mem[83][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19523_ (.CLK(clknet_leaf_48_clk),
    .D(_00821_),
    .Q(\cur_mb_mem[83][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19524_ (.CLK(clknet_leaf_52_clk),
    .D(_00822_),
    .Q(\cur_mb_mem[83][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19525_ (.CLK(clknet_leaf_63_clk),
    .D(_00823_),
    .Q(\cur_mb_mem[84][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19526_ (.CLK(clknet_leaf_130_clk),
    .D(_00824_),
    .Q(\cur_mb_mem[84][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19527_ (.CLK(clknet_leaf_68_clk),
    .D(_00825_),
    .Q(\cur_mb_mem[84][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19528_ (.CLK(clknet_leaf_96_clk),
    .D(_00826_),
    .Q(\cur_mb_mem[84][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19529_ (.CLK(clknet_leaf_99_clk),
    .D(_00827_),
    .Q(\cur_mb_mem[84][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19530_ (.CLK(clknet_leaf_99_clk),
    .D(_00828_),
    .Q(\cur_mb_mem[84][5] ));
 sky130_fd_sc_hd__dfxtp_2 _19531_ (.CLK(clknet_leaf_146_clk),
    .D(_00829_),
    .Q(\cur_mb_mem[84][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19532_ (.CLK(clknet_leaf_145_clk),
    .D(_00830_),
    .Q(\cur_mb_mem[84][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19533_ (.CLK(clknet_leaf_91_clk),
    .D(_00831_),
    .Q(\cur_mb_mem[85][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19534_ (.CLK(clknet_leaf_50_clk),
    .D(_00832_),
    .Q(\cur_mb_mem[85][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19535_ (.CLK(clknet_leaf_84_clk),
    .D(_00833_),
    .Q(\cur_mb_mem[85][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19536_ (.CLK(clknet_leaf_62_clk),
    .D(_00834_),
    .Q(\cur_mb_mem[85][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19537_ (.CLK(clknet_leaf_77_clk),
    .D(_00835_),
    .Q(\cur_mb_mem[85][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19538_ (.CLK(clknet_leaf_78_clk),
    .D(_00836_),
    .Q(\cur_mb_mem[85][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19539_ (.CLK(clknet_leaf_150_clk),
    .D(_00837_),
    .Q(\cur_mb_mem[85][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19540_ (.CLK(clknet_leaf_52_clk),
    .D(_00838_),
    .Q(\cur_mb_mem[85][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19541_ (.CLK(clknet_leaf_111_clk),
    .D(_00839_),
    .Q(\cur_mb_mem[86][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19542_ (.CLK(clknet_leaf_153_clk),
    .D(_00840_),
    .Q(\cur_mb_mem[86][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19543_ (.CLK(clknet_leaf_143_clk),
    .D(_00841_),
    .Q(\cur_mb_mem[86][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19544_ (.CLK(clknet_leaf_111_clk),
    .D(_00842_),
    .Q(\cur_mb_mem[86][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19545_ (.CLK(clknet_leaf_125_clk),
    .D(_00843_),
    .Q(\cur_mb_mem[86][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19546_ (.CLK(clknet_leaf_126_clk),
    .D(_00844_),
    .Q(\cur_mb_mem[86][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19547_ (.CLK(clknet_leaf_50_clk),
    .D(_00845_),
    .Q(\cur_mb_mem[86][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19548_ (.CLK(clknet_leaf_242_clk),
    .D(_00846_),
    .Q(\cur_mb_mem[86][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19549_ (.CLK(clknet_leaf_251_clk),
    .D(_00847_),
    .Q(\cur_mb_mem[87][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19550_ (.CLK(clknet_leaf_323_clk),
    .D(_00848_),
    .Q(\cur_mb_mem[87][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19551_ (.CLK(clknet_leaf_251_clk),
    .D(_00849_),
    .Q(\cur_mb_mem[87][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19552_ (.CLK(clknet_leaf_246_clk),
    .D(_00850_),
    .Q(\cur_mb_mem[87][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19553_ (.CLK(clknet_leaf_132_clk),
    .D(_00851_),
    .Q(\cur_mb_mem[87][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19554_ (.CLK(clknet_leaf_132_clk),
    .D(_00852_),
    .Q(\cur_mb_mem[87][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19555_ (.CLK(clknet_leaf_322_clk),
    .D(_00853_),
    .Q(\cur_mb_mem[87][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19556_ (.CLK(clknet_leaf_322_clk),
    .D(_00854_),
    .Q(\cur_mb_mem[87][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19557_ (.CLK(clknet_leaf_96_clk),
    .D(_00855_),
    .Q(\cur_mb_mem[88][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19558_ (.CLK(clknet_leaf_131_clk),
    .D(_00856_),
    .Q(\cur_mb_mem[88][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19559_ (.CLK(clknet_leaf_94_clk),
    .D(_00857_),
    .Q(\cur_mb_mem[88][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19560_ (.CLK(clknet_leaf_96_clk),
    .D(_00858_),
    .Q(\cur_mb_mem[88][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19561_ (.CLK(clknet_leaf_110_clk),
    .D(_00859_),
    .Q(\cur_mb_mem[88][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19562_ (.CLK(clknet_leaf_136_clk),
    .D(_00860_),
    .Q(\cur_mb_mem[88][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19563_ (.CLK(clknet_leaf_145_clk),
    .D(_00861_),
    .Q(\cur_mb_mem[88][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19564_ (.CLK(clknet_leaf_159_clk),
    .D(_00862_),
    .Q(\cur_mb_mem[88][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19565_ (.CLK(clknet_leaf_70_clk),
    .D(_00863_),
    .Q(\cur_mb_mem[89][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19566_ (.CLK(clknet_leaf_59_clk),
    .D(_00864_),
    .Q(\cur_mb_mem[89][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19567_ (.CLK(clknet_leaf_46_clk),
    .D(_00865_),
    .Q(\cur_mb_mem[89][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19568_ (.CLK(clknet_leaf_30_clk),
    .D(_00866_),
    .Q(\cur_mb_mem[89][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19569_ (.CLK(clknet_leaf_44_clk),
    .D(_00867_),
    .Q(\cur_mb_mem[89][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19570_ (.CLK(clknet_leaf_58_clk),
    .D(_00868_),
    .Q(\cur_mb_mem[89][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19571_ (.CLK(clknet_leaf_331_clk),
    .D(_00869_),
    .Q(\cur_mb_mem[89][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19572_ (.CLK(clknet_leaf_151_clk),
    .D(_00870_),
    .Q(\cur_mb_mem[89][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19573_ (.CLK(clknet_leaf_89_clk),
    .D(_00871_),
    .Q(\cur_mb_mem[90][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19574_ (.CLK(clknet_leaf_322_clk),
    .D(_00872_),
    .Q(\cur_mb_mem[90][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19575_ (.CLK(clknet_leaf_89_clk),
    .D(_00873_),
    .Q(\cur_mb_mem[90][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19576_ (.CLK(clknet_leaf_93_clk),
    .D(_00874_),
    .Q(\cur_mb_mem[90][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19577_ (.CLK(clknet_leaf_98_clk),
    .D(_00875_),
    .Q(\cur_mb_mem[90][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19578_ (.CLK(clknet_leaf_98_clk),
    .D(_00876_),
    .Q(\cur_mb_mem[90][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19579_ (.CLK(clknet_leaf_339_clk),
    .D(_00877_),
    .Q(\cur_mb_mem[90][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19580_ (.CLK(clknet_leaf_331_clk),
    .D(_00878_),
    .Q(\cur_mb_mem[90][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19581_ (.CLK(clknet_leaf_33_clk),
    .D(_00879_),
    .Q(\cur_mb_mem[91][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19582_ (.CLK(clknet_leaf_240_clk),
    .D(_00880_),
    .Q(\cur_mb_mem[91][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19583_ (.CLK(clknet_leaf_31_clk),
    .D(_00881_),
    .Q(\cur_mb_mem[91][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19584_ (.CLK(clknet_leaf_29_clk),
    .D(_00882_),
    .Q(\cur_mb_mem[91][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19585_ (.CLK(clknet_leaf_106_clk),
    .D(_00883_),
    .Q(\cur_mb_mem[91][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19586_ (.CLK(clknet_leaf_108_clk),
    .D(_00884_),
    .Q(\cur_mb_mem[91][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19587_ (.CLK(clknet_leaf_146_clk),
    .D(_00885_),
    .Q(\cur_mb_mem[91][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19588_ (.CLK(clknet_leaf_240_clk),
    .D(_00886_),
    .Q(\cur_mb_mem[91][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19589_ (.CLK(clknet_leaf_148_clk),
    .D(_00887_),
    .Q(\cur_mb_mem[92][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19590_ (.CLK(clknet_leaf_44_clk),
    .D(_00888_),
    .Q(\cur_mb_mem[92][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19591_ (.CLK(clknet_leaf_157_clk),
    .D(_00889_),
    .Q(\cur_mb_mem[92][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19592_ (.CLK(clknet_leaf_61_clk),
    .D(_00890_),
    .Q(\cur_mb_mem[92][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19593_ (.CLK(clknet_leaf_106_clk),
    .D(_00891_),
    .Q(\cur_mb_mem[92][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19594_ (.CLK(clknet_leaf_106_clk),
    .D(_00892_),
    .Q(\cur_mb_mem[92][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19595_ (.CLK(clknet_leaf_330_clk),
    .D(_00893_),
    .Q(\cur_mb_mem[92][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19596_ (.CLK(clknet_leaf_150_clk),
    .D(_00894_),
    .Q(\cur_mb_mem[92][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19597_ (.CLK(clknet_leaf_7_clk),
    .D(_00895_),
    .Q(\cur_mb_mem[93][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19598_ (.CLK(clknet_leaf_339_clk),
    .D(_00896_),
    .Q(\cur_mb_mem[93][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19599_ (.CLK(clknet_leaf_7_clk),
    .D(_00897_),
    .Q(\cur_mb_mem[93][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19600_ (.CLK(clknet_leaf_37_clk),
    .D(_00898_),
    .Q(\cur_mb_mem[93][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19601_ (.CLK(clknet_leaf_125_clk),
    .D(_00899_),
    .Q(\cur_mb_mem[93][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19602_ (.CLK(clknet_leaf_125_clk),
    .D(_00900_),
    .Q(\cur_mb_mem[93][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19603_ (.CLK(clknet_leaf_331_clk),
    .D(_00901_),
    .Q(\cur_mb_mem[93][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19604_ (.CLK(clknet_leaf_150_clk),
    .D(_00902_),
    .Q(\cur_mb_mem[93][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19605_ (.CLK(clknet_leaf_321_clk),
    .D(_00903_),
    .Q(\cur_mb_mem[94][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19606_ (.CLK(clknet_leaf_59_clk),
    .D(_00904_),
    .Q(\cur_mb_mem[94][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19607_ (.CLK(clknet_leaf_321_clk),
    .D(_00905_),
    .Q(\cur_mb_mem[94][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19608_ (.CLK(clknet_leaf_322_clk),
    .D(_00906_),
    .Q(\cur_mb_mem[94][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19609_ (.CLK(clknet_leaf_107_clk),
    .D(_00907_),
    .Q(\cur_mb_mem[94][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19610_ (.CLK(clknet_leaf_107_clk),
    .D(_00908_),
    .Q(\cur_mb_mem[94][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19611_ (.CLK(clknet_leaf_339_clk),
    .D(_00909_),
    .Q(\cur_mb_mem[94][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19612_ (.CLK(clknet_leaf_155_clk),
    .D(_00910_),
    .Q(\cur_mb_mem[94][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19613_ (.CLK(clknet_leaf_164_clk),
    .D(_00911_),
    .Q(\cur_mb_mem[95][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19614_ (.CLK(clknet_leaf_153_clk),
    .D(_00912_),
    .Q(\cur_mb_mem[95][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19615_ (.CLK(clknet_leaf_164_clk),
    .D(_00913_),
    .Q(\cur_mb_mem[95][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19616_ (.CLK(clknet_leaf_164_clk),
    .D(_00914_),
    .Q(\cur_mb_mem[95][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19617_ (.CLK(clknet_leaf_68_clk),
    .D(_00915_),
    .Q(\cur_mb_mem[95][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19618_ (.CLK(clknet_leaf_75_clk),
    .D(_00916_),
    .Q(\cur_mb_mem[95][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19619_ (.CLK(clknet_leaf_151_clk),
    .D(_00917_),
    .Q(\cur_mb_mem[95][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19620_ (.CLK(clknet_leaf_156_clk),
    .D(_00918_),
    .Q(\cur_mb_mem[95][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19621_ (.CLK(clknet_leaf_79_clk),
    .D(_00919_),
    .Q(\cur_mb_mem[96][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19622_ (.CLK(clknet_leaf_77_clk),
    .D(_00920_),
    .Q(\cur_mb_mem[96][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19623_ (.CLK(clknet_leaf_81_clk),
    .D(_00921_),
    .Q(\cur_mb_mem[96][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19624_ (.CLK(clknet_leaf_83_clk),
    .D(_00922_),
    .Q(\cur_mb_mem[96][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19625_ (.CLK(clknet_leaf_24_clk),
    .D(_00923_),
    .Q(\cur_mb_mem[96][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19626_ (.CLK(clknet_leaf_24_clk),
    .D(_00924_),
    .Q(\cur_mb_mem[96][5] ));
 sky130_fd_sc_hd__dfxtp_2 _19627_ (.CLK(clknet_leaf_83_clk),
    .D(_00925_),
    .Q(\cur_mb_mem[96][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19628_ (.CLK(clknet_leaf_83_clk),
    .D(_00926_),
    .Q(\cur_mb_mem[96][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19629_ (.CLK(clknet_leaf_83_clk),
    .D(_00927_),
    .Q(\cur_mb_mem[97][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19630_ (.CLK(clknet_leaf_82_clk),
    .D(_00928_),
    .Q(\cur_mb_mem[97][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19631_ (.CLK(clknet_leaf_80_clk),
    .D(_00929_),
    .Q(\cur_mb_mem[97][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19632_ (.CLK(clknet_leaf_81_clk),
    .D(_00930_),
    .Q(\cur_mb_mem[97][3] ));
 sky130_fd_sc_hd__dfxtp_2 _19633_ (.CLK(clknet_leaf_82_clk),
    .D(_00931_),
    .Q(\cur_mb_mem[97][4] ));
 sky130_fd_sc_hd__dfxtp_2 _19634_ (.CLK(clknet_leaf_80_clk),
    .D(_00932_),
    .Q(\cur_mb_mem[97][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19635_ (.CLK(clknet_leaf_21_clk),
    .D(_00933_),
    .Q(\cur_mb_mem[97][6] ));
 sky130_fd_sc_hd__dfxtp_4 _19636_ (.CLK(clknet_leaf_82_clk),
    .D(_00934_),
    .Q(\cur_mb_mem[97][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19637_ (.CLK(clknet_leaf_21_clk),
    .D(_00935_),
    .Q(\cur_mb_mem[98][0] ));
 sky130_fd_sc_hd__dfxtp_2 _19638_ (.CLK(clknet_leaf_23_clk),
    .D(_00936_),
    .Q(\cur_mb_mem[98][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19639_ (.CLK(clknet_leaf_21_clk),
    .D(_00937_),
    .Q(\cur_mb_mem[98][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19640_ (.CLK(clknet_leaf_23_clk),
    .D(_00938_),
    .Q(\cur_mb_mem[98][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19641_ (.CLK(clknet_leaf_82_clk),
    .D(_00939_),
    .Q(\cur_mb_mem[98][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19642_ (.CLK(clknet_leaf_79_clk),
    .D(_00940_),
    .Q(\cur_mb_mem[98][5] ));
 sky130_fd_sc_hd__dfxtp_2 _19643_ (.CLK(clknet_leaf_86_clk),
    .D(_00941_),
    .Q(\cur_mb_mem[98][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19644_ (.CLK(clknet_leaf_17_clk),
    .D(_00942_),
    .Q(\cur_mb_mem[98][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19645_ (.CLK(clknet_leaf_317_clk),
    .D(_00943_),
    .Q(\cur_mb_mem[99][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19646_ (.CLK(clknet_leaf_342_clk),
    .D(_00944_),
    .Q(\cur_mb_mem[99][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19647_ (.CLK(clknet_leaf_317_clk),
    .D(_00945_),
    .Q(\cur_mb_mem[99][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19648_ (.CLK(clknet_leaf_317_clk),
    .D(_00946_),
    .Q(\cur_mb_mem[99][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19649_ (.CLK(clknet_leaf_75_clk),
    .D(_00947_),
    .Q(\cur_mb_mem[99][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19650_ (.CLK(clknet_leaf_75_clk),
    .D(_00948_),
    .Q(\cur_mb_mem[99][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19651_ (.CLK(clknet_leaf_324_clk),
    .D(_00949_),
    .Q(\cur_mb_mem[99][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19652_ (.CLK(clknet_leaf_319_clk),
    .D(_00950_),
    .Q(\cur_mb_mem[99][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19653_ (.CLK(clknet_leaf_85_clk),
    .D(_00951_),
    .Q(\cur_mb_mem[100][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19654_ (.CLK(clknet_leaf_81_clk),
    .D(_00952_),
    .Q(\cur_mb_mem[100][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19655_ (.CLK(clknet_leaf_86_clk),
    .D(_00953_),
    .Q(\cur_mb_mem[100][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19656_ (.CLK(clknet_leaf_85_clk),
    .D(_00954_),
    .Q(\cur_mb_mem[100][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19657_ (.CLK(clknet_leaf_23_clk),
    .D(_00955_),
    .Q(\cur_mb_mem[100][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19658_ (.CLK(clknet_leaf_79_clk),
    .D(_00956_),
    .Q(\cur_mb_mem[100][5] ));
 sky130_fd_sc_hd__dfxtp_2 _19659_ (.CLK(clknet_leaf_86_clk),
    .D(_00957_),
    .Q(\cur_mb_mem[100][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19660_ (.CLK(clknet_leaf_85_clk),
    .D(_00958_),
    .Q(\cur_mb_mem[100][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19661_ (.CLK(clknet_leaf_166_clk),
    .D(_00959_),
    .Q(\cur_mb_mem[101][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19662_ (.CLK(clknet_leaf_323_clk),
    .D(_00960_),
    .Q(\cur_mb_mem[101][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19663_ (.CLK(clknet_leaf_166_clk),
    .D(_00961_),
    .Q(\cur_mb_mem[101][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19664_ (.CLK(clknet_leaf_166_clk),
    .D(_00962_),
    .Q(\cur_mb_mem[101][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19665_ (.CLK(clknet_leaf_29_clk),
    .D(_00963_),
    .Q(\cur_mb_mem[101][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19666_ (.CLK(clknet_leaf_27_clk),
    .D(_00964_),
    .Q(\cur_mb_mem[101][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19667_ (.CLK(clknet_leaf_146_clk),
    .D(_00965_),
    .Q(\cur_mb_mem[101][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19668_ (.CLK(clknet_leaf_154_clk),
    .D(_00966_),
    .Q(\cur_mb_mem[101][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19669_ (.CLK(clknet_leaf_74_clk),
    .D(_00967_),
    .Q(\cur_mb_mem[102][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19670_ (.CLK(clknet_leaf_40_clk),
    .D(_00968_),
    .Q(\cur_mb_mem[102][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19671_ (.CLK(clknet_leaf_74_clk),
    .D(_00969_),
    .Q(\cur_mb_mem[102][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19672_ (.CLK(clknet_leaf_75_clk),
    .D(_00970_),
    .Q(\cur_mb_mem[102][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19673_ (.CLK(clknet_leaf_75_clk),
    .D(_00971_),
    .Q(\cur_mb_mem[102][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19674_ (.CLK(clknet_leaf_74_clk),
    .D(_00972_),
    .Q(\cur_mb_mem[102][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19675_ (.CLK(clknet_leaf_343_clk),
    .D(_00973_),
    .Q(\cur_mb_mem[102][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19676_ (.CLK(clknet_leaf_343_clk),
    .D(_00974_),
    .Q(\cur_mb_mem[102][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19677_ (.CLK(clknet_leaf_93_clk),
    .D(_00975_),
    .Q(\cur_mb_mem[103][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19678_ (.CLK(clknet_leaf_157_clk),
    .D(_00976_),
    .Q(\cur_mb_mem[103][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19679_ (.CLK(clknet_leaf_64_clk),
    .D(_00977_),
    .Q(\cur_mb_mem[103][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19680_ (.CLK(clknet_leaf_89_clk),
    .D(_00978_),
    .Q(\cur_mb_mem[103][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19681_ (.CLK(clknet_leaf_84_clk),
    .D(_00979_),
    .Q(\cur_mb_mem[103][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19682_ (.CLK(clknet_leaf_76_clk),
    .D(_00980_),
    .Q(\cur_mb_mem[103][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19683_ (.CLK(clknet_leaf_320_clk),
    .D(_00981_),
    .Q(\cur_mb_mem[103][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19684_ (.CLK(clknet_leaf_327_clk),
    .D(_00982_),
    .Q(\cur_mb_mem[103][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19685_ (.CLK(clknet_leaf_86_clk),
    .D(_00983_),
    .Q(\cur_mb_mem[104][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19686_ (.CLK(clknet_leaf_80_clk),
    .D(_00984_),
    .Q(\cur_mb_mem[104][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19687_ (.CLK(clknet_leaf_86_clk),
    .D(_00985_),
    .Q(\cur_mb_mem[104][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19688_ (.CLK(clknet_leaf_86_clk),
    .D(_00986_),
    .Q(\cur_mb_mem[104][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19689_ (.CLK(clknet_leaf_394_clk),
    .D(_00987_),
    .Q(\cur_mb_mem[104][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19690_ (.CLK(clknet_leaf_394_clk),
    .D(_00988_),
    .Q(\cur_mb_mem[104][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19691_ (.CLK(clknet_leaf_21_clk),
    .D(_00989_),
    .Q(\cur_mb_mem[104][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19692_ (.CLK(clknet_leaf_21_clk),
    .D(_00990_),
    .Q(\cur_mb_mem[104][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19693_ (.CLK(clknet_leaf_67_clk),
    .D(_00991_),
    .Q(\cur_mb_mem[105][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19694_ (.CLK(clknet_leaf_346_clk),
    .D(_00992_),
    .Q(\cur_mb_mem[105][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19695_ (.CLK(clknet_leaf_140_clk),
    .D(_00993_),
    .Q(\cur_mb_mem[105][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19696_ (.CLK(clknet_leaf_65_clk),
    .D(_00994_),
    .Q(\cur_mb_mem[105][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19697_ (.CLK(clknet_leaf_28_clk),
    .D(_00995_),
    .Q(\cur_mb_mem[105][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19698_ (.CLK(clknet_leaf_28_clk),
    .D(_00996_),
    .Q(\cur_mb_mem[105][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19699_ (.CLK(clknet_leaf_158_clk),
    .D(_00997_),
    .Q(\cur_mb_mem[105][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19700_ (.CLK(clknet_leaf_342_clk),
    .D(_00998_),
    .Q(\cur_mb_mem[105][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19701_ (.CLK(clknet_leaf_91_clk),
    .D(_00999_),
    .Q(\cur_mb_mem[106][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19702_ (.CLK(clknet_leaf_29_clk),
    .D(_01000_),
    .Q(\cur_mb_mem[106][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19703_ (.CLK(clknet_leaf_140_clk),
    .D(_01001_),
    .Q(\cur_mb_mem[106][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19704_ (.CLK(clknet_leaf_65_clk),
    .D(_01002_),
    .Q(\cur_mb_mem[106][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19705_ (.CLK(clknet_leaf_76_clk),
    .D(_01003_),
    .Q(\cur_mb_mem[106][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19706_ (.CLK(clknet_leaf_74_clk),
    .D(_01004_),
    .Q(\cur_mb_mem[106][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19707_ (.CLK(clknet_leaf_142_clk),
    .D(_01005_),
    .Q(\cur_mb_mem[106][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19708_ (.CLK(clknet_leaf_141_clk),
    .D(_01006_),
    .Q(\cur_mb_mem[106][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19709_ (.CLK(clknet_leaf_9_clk),
    .D(_01007_),
    .Q(\cur_mb_mem[107][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19710_ (.CLK(clknet_leaf_72_clk),
    .D(_01008_),
    .Q(\cur_mb_mem[107][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19711_ (.CLK(clknet_leaf_13_clk),
    .D(_01009_),
    .Q(\cur_mb_mem[107][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19712_ (.CLK(clknet_leaf_26_clk),
    .D(_01010_),
    .Q(\cur_mb_mem[107][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19713_ (.CLK(clknet_leaf_62_clk),
    .D(_01011_),
    .Q(\cur_mb_mem[107][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19714_ (.CLK(clknet_leaf_62_clk),
    .D(_01012_),
    .Q(\cur_mb_mem[107][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19715_ (.CLK(clknet_leaf_148_clk),
    .D(_01013_),
    .Q(\cur_mb_mem[107][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19716_ (.CLK(clknet_leaf_53_clk),
    .D(_01014_),
    .Q(\cur_mb_mem[107][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19717_ (.CLK(clknet_leaf_87_clk),
    .D(_01015_),
    .Q(\cur_mb_mem[108][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19718_ (.CLK(clknet_leaf_62_clk),
    .D(_01016_),
    .Q(\cur_mb_mem[108][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19719_ (.CLK(clknet_leaf_87_clk),
    .D(_01017_),
    .Q(\cur_mb_mem[108][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19720_ (.CLK(clknet_leaf_88_clk),
    .D(_01018_),
    .Q(\cur_mb_mem[108][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19721_ (.CLK(clknet_leaf_377_clk),
    .D(_01019_),
    .Q(\cur_mb_mem[108][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19722_ (.CLK(clknet_leaf_374_clk),
    .D(_01020_),
    .Q(\cur_mb_mem[108][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19723_ (.CLK(clknet_leaf_159_clk),
    .D(_01021_),
    .Q(\cur_mb_mem[108][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19724_ (.CLK(clknet_leaf_359_clk),
    .D(_01022_),
    .Q(\cur_mb_mem[108][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19725_ (.CLK(clknet_leaf_29_clk),
    .D(_01023_),
    .Q(\cur_mb_mem[109][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19726_ (.CLK(clknet_leaf_60_clk),
    .D(_01024_),
    .Q(\cur_mb_mem[109][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19727_ (.CLK(clknet_leaf_73_clk),
    .D(_01025_),
    .Q(\cur_mb_mem[109][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19728_ (.CLK(clknet_leaf_69_clk),
    .D(_01026_),
    .Q(\cur_mb_mem[109][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19729_ (.CLK(clknet_leaf_58_clk),
    .D(_01027_),
    .Q(\cur_mb_mem[109][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19730_ (.CLK(clknet_leaf_57_clk),
    .D(_01028_),
    .Q(\cur_mb_mem[109][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19731_ (.CLK(clknet_leaf_70_clk),
    .D(_01029_),
    .Q(\cur_mb_mem[109][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19732_ (.CLK(clknet_leaf_147_clk),
    .D(_01030_),
    .Q(\cur_mb_mem[109][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19733_ (.CLK(clknet_leaf_29_clk),
    .D(_01031_),
    .Q(\cur_mb_mem[110][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19734_ (.CLK(clknet_leaf_49_clk),
    .D(_01032_),
    .Q(\cur_mb_mem[110][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19735_ (.CLK(clknet_leaf_73_clk),
    .D(_01033_),
    .Q(\cur_mb_mem[110][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19736_ (.CLK(clknet_leaf_69_clk),
    .D(_01034_),
    .Q(\cur_mb_mem[110][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19737_ (.CLK(clknet_leaf_58_clk),
    .D(_01035_),
    .Q(\cur_mb_mem[110][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19738_ (.CLK(clknet_leaf_57_clk),
    .D(_01036_),
    .Q(\cur_mb_mem[110][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19739_ (.CLK(clknet_leaf_29_clk),
    .D(_01037_),
    .Q(\cur_mb_mem[110][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19740_ (.CLK(clknet_leaf_149_clk),
    .D(_01038_),
    .Q(\cur_mb_mem[110][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19741_ (.CLK(clknet_leaf_93_clk),
    .D(_01039_),
    .Q(\cur_mb_mem[111][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19742_ (.CLK(clknet_leaf_307_clk),
    .D(_01040_),
    .Q(\cur_mb_mem[111][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19743_ (.CLK(clknet_leaf_64_clk),
    .D(_01041_),
    .Q(\cur_mb_mem[111][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19744_ (.CLK(clknet_leaf_92_clk),
    .D(_01042_),
    .Q(\cur_mb_mem[111][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19745_ (.CLK(clknet_leaf_385_clk),
    .D(_01043_),
    .Q(\cur_mb_mem[111][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19746_ (.CLK(clknet_leaf_385_clk),
    .D(_01044_),
    .Q(\cur_mb_mem[111][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19747_ (.CLK(clknet_leaf_305_clk),
    .D(_01045_),
    .Q(\cur_mb_mem[111][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19748_ (.CLK(clknet_leaf_301_clk),
    .D(_01046_),
    .Q(\cur_mb_mem[111][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19749_ (.CLK(clknet_leaf_81_clk),
    .D(_01047_),
    .Q(\cur_mb_mem[112][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19750_ (.CLK(clknet_leaf_78_clk),
    .D(_01048_),
    .Q(\cur_mb_mem[112][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19751_ (.CLK(clknet_leaf_79_clk),
    .D(_01049_),
    .Q(\cur_mb_mem[112][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19752_ (.CLK(clknet_leaf_81_clk),
    .D(_01050_),
    .Q(\cur_mb_mem[112][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19753_ (.CLK(clknet_leaf_20_clk),
    .D(_01051_),
    .Q(\cur_mb_mem[112][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19754_ (.CLK(clknet_leaf_20_clk),
    .D(_01052_),
    .Q(\cur_mb_mem[112][5] ));
 sky130_fd_sc_hd__dfxtp_2 _19755_ (.CLK(clknet_leaf_22_clk),
    .D(_01053_),
    .Q(\cur_mb_mem[112][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19756_ (.CLK(clknet_leaf_17_clk),
    .D(_01054_),
    .Q(\cur_mb_mem[112][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19757_ (.CLK(clknet_leaf_22_clk),
    .D(_01055_),
    .Q(\cur_mb_mem[113][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19758_ (.CLK(clknet_leaf_23_clk),
    .D(_01056_),
    .Q(\cur_mb_mem[113][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19759_ (.CLK(clknet_leaf_24_clk),
    .D(_01057_),
    .Q(\cur_mb_mem[113][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19760_ (.CLK(clknet_leaf_22_clk),
    .D(_01058_),
    .Q(\cur_mb_mem[113][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19761_ (.CLK(clknet_leaf_16_clk),
    .D(_01059_),
    .Q(\cur_mb_mem[113][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19762_ (.CLK(clknet_leaf_16_clk),
    .D(_01060_),
    .Q(\cur_mb_mem[113][5] ));
 sky130_fd_sc_hd__dfxtp_2 _19763_ (.CLK(clknet_leaf_24_clk),
    .D(_01061_),
    .Q(\cur_mb_mem[113][6] ));
 sky130_fd_sc_hd__dfxtp_4 _19764_ (.CLK(clknet_leaf_21_clk),
    .D(_01062_),
    .Q(\cur_mb_mem[113][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19765_ (.CLK(clknet_leaf_23_clk),
    .D(_01063_),
    .Q(\cur_mb_mem[114][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19766_ (.CLK(clknet_leaf_23_clk),
    .D(_01064_),
    .Q(\cur_mb_mem[114][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19767_ (.CLK(clknet_leaf_79_clk),
    .D(_01065_),
    .Q(\cur_mb_mem[114][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19768_ (.CLK(clknet_leaf_80_clk),
    .D(_01066_),
    .Q(\cur_mb_mem[114][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19769_ (.CLK(clknet_leaf_16_clk),
    .D(_01067_),
    .Q(\cur_mb_mem[114][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19770_ (.CLK(clknet_leaf_16_clk),
    .D(_01068_),
    .Q(\cur_mb_mem[114][5] ));
 sky130_fd_sc_hd__dfxtp_2 _19771_ (.CLK(clknet_leaf_79_clk),
    .D(_01069_),
    .Q(\cur_mb_mem[114][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19772_ (.CLK(clknet_leaf_82_clk),
    .D(_01070_),
    .Q(\cur_mb_mem[114][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19773_ (.CLK(clknet_leaf_87_clk),
    .D(_01071_),
    .Q(\cur_mb_mem[115][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19774_ (.CLK(clknet_leaf_36_clk),
    .D(_01072_),
    .Q(\cur_mb_mem[115][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19775_ (.CLK(clknet_leaf_87_clk),
    .D(_01073_),
    .Q(\cur_mb_mem[115][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19776_ (.CLK(clknet_leaf_91_clk),
    .D(_01074_),
    .Q(\cur_mb_mem[115][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19777_ (.CLK(clknet_leaf_13_clk),
    .D(_01075_),
    .Q(\cur_mb_mem[115][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19778_ (.CLK(clknet_leaf_0_clk),
    .D(_01076_),
    .Q(\cur_mb_mem[115][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19779_ (.CLK(clknet_leaf_13_clk),
    .D(_01077_),
    .Q(\cur_mb_mem[115][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19780_ (.CLK(clknet_leaf_345_clk),
    .D(_01078_),
    .Q(\cur_mb_mem[115][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19781_ (.CLK(clknet_leaf_22_clk),
    .D(_01079_),
    .Q(\cur_mb_mem[116][0] ));
 sky130_fd_sc_hd__dfxtp_2 _19782_ (.CLK(clknet_leaf_80_clk),
    .D(_01080_),
    .Q(\cur_mb_mem[116][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19783_ (.CLK(clknet_leaf_21_clk),
    .D(_01081_),
    .Q(\cur_mb_mem[116][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19784_ (.CLK(clknet_leaf_22_clk),
    .D(_01082_),
    .Q(\cur_mb_mem[116][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19785_ (.CLK(clknet_leaf_21_clk),
    .D(_01083_),
    .Q(\cur_mb_mem[116][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19786_ (.CLK(clknet_leaf_22_clk),
    .D(_01084_),
    .Q(\cur_mb_mem[116][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19787_ (.CLK(clknet_leaf_79_clk),
    .D(_01085_),
    .Q(\cur_mb_mem[116][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19788_ (.CLK(clknet_leaf_86_clk),
    .D(_01086_),
    .Q(\cur_mb_mem[116][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19789_ (.CLK(clknet_leaf_76_clk),
    .D(_01087_),
    .Q(\cur_mb_mem[117][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19790_ (.CLK(clknet_leaf_16_clk),
    .D(_01088_),
    .Q(\cur_mb_mem[117][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19791_ (.CLK(clknet_leaf_78_clk),
    .D(_01089_),
    .Q(\cur_mb_mem[117][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19792_ (.CLK(clknet_leaf_76_clk),
    .D(_01090_),
    .Q(\cur_mb_mem[117][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19793_ (.CLK(clknet_leaf_17_clk),
    .D(_01091_),
    .Q(\cur_mb_mem[117][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19794_ (.CLK(clknet_leaf_17_clk),
    .D(_01092_),
    .Q(\cur_mb_mem[117][5] ));
 sky130_fd_sc_hd__dfxtp_2 _19795_ (.CLK(clknet_leaf_17_clk),
    .D(_01093_),
    .Q(\cur_mb_mem[117][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19796_ (.CLK(clknet_leaf_34_clk),
    .D(_01094_),
    .Q(\cur_mb_mem[117][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19797_ (.CLK(clknet_leaf_308_clk),
    .D(_01095_),
    .Q(\cur_mb_mem[118][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19798_ (.CLK(clknet_leaf_333_clk),
    .D(_01096_),
    .Q(\cur_mb_mem[118][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19799_ (.CLK(clknet_leaf_309_clk),
    .D(_01097_),
    .Q(\cur_mb_mem[118][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19800_ (.CLK(clknet_leaf_307_clk),
    .D(_01098_),
    .Q(\cur_mb_mem[118][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19801_ (.CLK(clknet_leaf_17_clk),
    .D(_01099_),
    .Q(\cur_mb_mem[118][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19802_ (.CLK(clknet_leaf_17_clk),
    .D(_01100_),
    .Q(\cur_mb_mem[118][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19803_ (.CLK(clknet_leaf_393_clk),
    .D(_01101_),
    .Q(\cur_mb_mem[118][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19804_ (.CLK(clknet_leaf_337_clk),
    .D(_01102_),
    .Q(\cur_mb_mem[118][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19805_ (.CLK(clknet_leaf_313_clk),
    .D(_01103_),
    .Q(\cur_mb_mem[119][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19806_ (.CLK(clknet_leaf_319_clk),
    .D(_01104_),
    .Q(\cur_mb_mem[119][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19807_ (.CLK(clknet_leaf_313_clk),
    .D(_01105_),
    .Q(\cur_mb_mem[119][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19808_ (.CLK(clknet_leaf_11_clk),
    .D(_01106_),
    .Q(\cur_mb_mem[119][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19809_ (.CLK(clknet_leaf_15_clk),
    .D(_01107_),
    .Q(\cur_mb_mem[119][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19810_ (.CLK(clknet_leaf_15_clk),
    .D(_01108_),
    .Q(\cur_mb_mem[119][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19811_ (.CLK(clknet_leaf_309_clk),
    .D(_01109_),
    .Q(\cur_mb_mem[119][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19812_ (.CLK(clknet_leaf_320_clk),
    .D(_01110_),
    .Q(\cur_mb_mem[119][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19813_ (.CLK(clknet_leaf_81_clk),
    .D(_01111_),
    .Q(\cur_mb_mem[120][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19814_ (.CLK(clknet_leaf_83_clk),
    .D(_01112_),
    .Q(\cur_mb_mem[120][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19815_ (.CLK(clknet_leaf_80_clk),
    .D(_01113_),
    .Q(\cur_mb_mem[120][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19816_ (.CLK(clknet_leaf_81_clk),
    .D(_01114_),
    .Q(\cur_mb_mem[120][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19817_ (.CLK(clknet_leaf_394_clk),
    .D(_01115_),
    .Q(\cur_mb_mem[120][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19818_ (.CLK(clknet_leaf_394_clk),
    .D(_01116_),
    .Q(\cur_mb_mem[120][5] ));
 sky130_fd_sc_hd__dfxtp_2 _19819_ (.CLK(clknet_leaf_81_clk),
    .D(_01117_),
    .Q(\cur_mb_mem[120][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19820_ (.CLK(clknet_leaf_21_clk),
    .D(_01118_),
    .Q(\cur_mb_mem[120][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19821_ (.CLK(clknet_leaf_83_clk),
    .D(_01119_),
    .Q(\cur_mb_mem[121][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19822_ (.CLK(clknet_leaf_19_clk),
    .D(_01120_),
    .Q(\cur_mb_mem[121][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19823_ (.CLK(clknet_leaf_84_clk),
    .D(_01121_),
    .Q(\cur_mb_mem[121][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19824_ (.CLK(clknet_leaf_91_clk),
    .D(_01122_),
    .Q(\cur_mb_mem[121][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19825_ (.CLK(clknet_leaf_20_clk),
    .D(_01123_),
    .Q(\cur_mb_mem[121][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19826_ (.CLK(clknet_leaf_19_clk),
    .D(_01124_),
    .Q(\cur_mb_mem[121][5] ));
 sky130_fd_sc_hd__dfxtp_2 _19827_ (.CLK(clknet_leaf_19_clk),
    .D(_01125_),
    .Q(\cur_mb_mem[121][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19828_ (.CLK(clknet_leaf_34_clk),
    .D(_01126_),
    .Q(\cur_mb_mem[121][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19829_ (.CLK(clknet_leaf_391_clk),
    .D(_01127_),
    .Q(\cur_mb_mem[122][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19830_ (.CLK(clknet_leaf_16_clk),
    .D(_01128_),
    .Q(\cur_mb_mem[122][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19831_ (.CLK(clknet_leaf_2_clk),
    .D(_01129_),
    .Q(\cur_mb_mem[122][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19832_ (.CLK(clknet_leaf_391_clk),
    .D(_01130_),
    .Q(\cur_mb_mem[122][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19833_ (.CLK(clknet_leaf_15_clk),
    .D(_01131_),
    .Q(\cur_mb_mem[122][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19834_ (.CLK(clknet_leaf_15_clk),
    .D(_01132_),
    .Q(\cur_mb_mem[122][5] ));
 sky130_fd_sc_hd__dfxtp_2 _19835_ (.CLK(clknet_leaf_393_clk),
    .D(_01133_),
    .Q(\cur_mb_mem[122][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19836_ (.CLK(clknet_leaf_10_clk),
    .D(_01134_),
    .Q(\cur_mb_mem[122][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19837_ (.CLK(clknet_leaf_8_clk),
    .D(_01135_),
    .Q(\cur_mb_mem[123][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19838_ (.CLK(clknet_leaf_32_clk),
    .D(_01136_),
    .Q(\cur_mb_mem[123][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19839_ (.CLK(clknet_leaf_9_clk),
    .D(_01137_),
    .Q(\cur_mb_mem[123][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19840_ (.CLK(clknet_leaf_8_clk),
    .D(_01138_),
    .Q(\cur_mb_mem[123][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19841_ (.CLK(clknet_leaf_19_clk),
    .D(_01139_),
    .Q(\cur_mb_mem[123][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19842_ (.CLK(clknet_leaf_18_clk),
    .D(_01140_),
    .Q(\cur_mb_mem[123][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19843_ (.CLK(clknet_leaf_17_clk),
    .D(_01141_),
    .Q(\cur_mb_mem[123][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19844_ (.CLK(clknet_leaf_36_clk),
    .D(_01142_),
    .Q(\cur_mb_mem[123][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19845_ (.CLK(clknet_leaf_3_clk),
    .D(_01143_),
    .Q(\cur_mb_mem[124][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19846_ (.CLK(clknet_leaf_15_clk),
    .D(_01144_),
    .Q(\cur_mb_mem[124][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19847_ (.CLK(clknet_leaf_392_clk),
    .D(_01145_),
    .Q(\cur_mb_mem[124][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19848_ (.CLK(clknet_leaf_392_clk),
    .D(_01146_),
    .Q(\cur_mb_mem[124][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19849_ (.CLK(clknet_leaf_392_clk),
    .D(_01147_),
    .Q(\cur_mb_mem[124][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19850_ (.CLK(clknet_leaf_393_clk),
    .D(_01148_),
    .Q(\cur_mb_mem[124][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19851_ (.CLK(clknet_leaf_394_clk),
    .D(_01149_),
    .Q(\cur_mb_mem[124][6] ));
 sky130_fd_sc_hd__dfxtp_2 _19852_ (.CLK(clknet_leaf_9_clk),
    .D(_01150_),
    .Q(\cur_mb_mem[124][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19853_ (.CLK(clknet_leaf_391_clk),
    .D(_01151_),
    .Q(\cur_mb_mem[125][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19854_ (.CLK(clknet_leaf_394_clk),
    .D(_01152_),
    .Q(\cur_mb_mem[125][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19855_ (.CLK(clknet_leaf_392_clk),
    .D(_01153_),
    .Q(\cur_mb_mem[125][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19856_ (.CLK(clknet_leaf_391_clk),
    .D(_01154_),
    .Q(\cur_mb_mem[125][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19857_ (.CLK(clknet_leaf_392_clk),
    .D(_01155_),
    .Q(\cur_mb_mem[125][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19858_ (.CLK(clknet_leaf_392_clk),
    .D(_01156_),
    .Q(\cur_mb_mem[125][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19859_ (.CLK(clknet_leaf_393_clk),
    .D(_01157_),
    .Q(\cur_mb_mem[125][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19860_ (.CLK(clknet_leaf_4_clk),
    .D(_01158_),
    .Q(\cur_mb_mem[125][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19861_ (.CLK(clknet_leaf_83_clk),
    .D(_01159_),
    .Q(\cur_mb_mem[126][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19862_ (.CLK(clknet_leaf_380_clk),
    .D(_01160_),
    .Q(\cur_mb_mem[126][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19863_ (.CLK(clknet_leaf_84_clk),
    .D(_01161_),
    .Q(\cur_mb_mem[126][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19864_ (.CLK(clknet_leaf_91_clk),
    .D(_01162_),
    .Q(\cur_mb_mem[126][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19865_ (.CLK(clknet_leaf_15_clk),
    .D(_01163_),
    .Q(\cur_mb_mem[126][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19866_ (.CLK(clknet_leaf_15_clk),
    .D(_01164_),
    .Q(\cur_mb_mem[126][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19867_ (.CLK(clknet_leaf_39_clk),
    .D(_01165_),
    .Q(\cur_mb_mem[126][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19868_ (.CLK(clknet_leaf_380_clk),
    .D(_01166_),
    .Q(\cur_mb_mem[126][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19869_ (.CLK(clknet_leaf_311_clk),
    .D(_01167_),
    .Q(\cur_mb_mem[127][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19870_ (.CLK(clknet_leaf_308_clk),
    .D(_01168_),
    .Q(\cur_mb_mem[127][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19871_ (.CLK(clknet_leaf_310_clk),
    .D(_01169_),
    .Q(\cur_mb_mem[127][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19872_ (.CLK(clknet_leaf_287_clk),
    .D(_01170_),
    .Q(\cur_mb_mem[127][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19873_ (.CLK(clknet_leaf_280_clk),
    .D(_01171_),
    .Q(\cur_mb_mem[127][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19874_ (.CLK(clknet_leaf_280_clk),
    .D(_01172_),
    .Q(\cur_mb_mem[127][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19875_ (.CLK(clknet_leaf_309_clk),
    .D(_01173_),
    .Q(\cur_mb_mem[127][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19876_ (.CLK(clknet_leaf_304_clk),
    .D(_01174_),
    .Q(\cur_mb_mem[127][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19877_ (.CLK(clknet_leaf_227_clk),
    .D(_01175_),
    .Q(\cur_mb_mem[128][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19878_ (.CLK(clknet_leaf_232_clk),
    .D(_01176_),
    .Q(\cur_mb_mem[128][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19879_ (.CLK(clknet_leaf_227_clk),
    .D(_01177_),
    .Q(\cur_mb_mem[128][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19880_ (.CLK(clknet_leaf_228_clk),
    .D(_01178_),
    .Q(\cur_mb_mem[128][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19881_ (.CLK(clknet_leaf_228_clk),
    .D(_01179_),
    .Q(\cur_mb_mem[128][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19882_ (.CLK(clknet_leaf_229_clk),
    .D(_01180_),
    .Q(\cur_mb_mem[128][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19883_ (.CLK(clknet_leaf_165_clk),
    .D(_01181_),
    .Q(\cur_mb_mem[128][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19884_ (.CLK(clknet_leaf_164_clk),
    .D(_01182_),
    .Q(\cur_mb_mem[128][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19885_ (.CLK(clknet_leaf_169_clk),
    .D(_01183_),
    .Q(\cur_mb_mem[129][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19886_ (.CLK(clknet_leaf_127_clk),
    .D(_01184_),
    .Q(\cur_mb_mem[129][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19887_ (.CLK(clknet_leaf_168_clk),
    .D(_01185_),
    .Q(\cur_mb_mem[129][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19888_ (.CLK(clknet_leaf_193_clk),
    .D(_01186_),
    .Q(\cur_mb_mem[129][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19889_ (.CLK(clknet_leaf_228_clk),
    .D(_01187_),
    .Q(\cur_mb_mem[129][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19890_ (.CLK(clknet_leaf_229_clk),
    .D(_01188_),
    .Q(\cur_mb_mem[129][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19891_ (.CLK(clknet_leaf_170_clk),
    .D(_01189_),
    .Q(\cur_mb_mem[129][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19892_ (.CLK(clknet_leaf_145_clk),
    .D(_01190_),
    .Q(\cur_mb_mem[129][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19893_ (.CLK(clknet_leaf_142_clk),
    .D(_01191_),
    .Q(\cur_mb_mem[130][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19894_ (.CLK(clknet_leaf_148_clk),
    .D(_01192_),
    .Q(\cur_mb_mem[130][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19895_ (.CLK(clknet_leaf_161_clk),
    .D(_01193_),
    .Q(\cur_mb_mem[130][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19896_ (.CLK(clknet_leaf_141_clk),
    .D(_01194_),
    .Q(\cur_mb_mem[130][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19897_ (.CLK(clknet_leaf_168_clk),
    .D(_01195_),
    .Q(\cur_mb_mem[130][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19898_ (.CLK(clknet_leaf_168_clk),
    .D(_01196_),
    .Q(\cur_mb_mem[130][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19899_ (.CLK(clknet_leaf_150_clk),
    .D(_01197_),
    .Q(\cur_mb_mem[130][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19900_ (.CLK(clknet_leaf_156_clk),
    .D(_01198_),
    .Q(\cur_mb_mem[130][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19901_ (.CLK(clknet_leaf_262_clk),
    .D(_01199_),
    .Q(\cur_mb_mem[131][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19902_ (.CLK(clknet_leaf_232_clk),
    .D(_01200_),
    .Q(\cur_mb_mem[131][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19903_ (.CLK(clknet_leaf_248_clk),
    .D(_01201_),
    .Q(\cur_mb_mem[131][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19904_ (.CLK(clknet_leaf_262_clk),
    .D(_01202_),
    .Q(\cur_mb_mem[131][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19905_ (.CLK(clknet_leaf_229_clk),
    .D(_01203_),
    .Q(\cur_mb_mem[131][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19906_ (.CLK(clknet_leaf_229_clk),
    .D(_01204_),
    .Q(\cur_mb_mem[131][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19907_ (.CLK(clknet_leaf_235_clk),
    .D(_01205_),
    .Q(\cur_mb_mem[131][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19908_ (.CLK(clknet_leaf_235_clk),
    .D(_01206_),
    .Q(\cur_mb_mem[131][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19909_ (.CLK(clknet_leaf_111_clk),
    .D(_01207_),
    .Q(\cur_mb_mem[132][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19910_ (.CLK(clknet_leaf_61_clk),
    .D(_01208_),
    .Q(\cur_mb_mem[132][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19911_ (.CLK(clknet_leaf_144_clk),
    .D(_01209_),
    .Q(\cur_mb_mem[132][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19912_ (.CLK(clknet_leaf_111_clk),
    .D(_01210_),
    .Q(\cur_mb_mem[132][3] ));
 sky130_fd_sc_hd__dfxtp_2 _19913_ (.CLK(clknet_leaf_85_clk),
    .D(_01211_),
    .Q(\cur_mb_mem[132][4] ));
 sky130_fd_sc_hd__dfxtp_2 _19914_ (.CLK(clknet_leaf_85_clk),
    .D(_01212_),
    .Q(\cur_mb_mem[132][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19915_ (.CLK(clknet_leaf_177_clk),
    .D(_01213_),
    .Q(\cur_mb_mem[132][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19916_ (.CLK(clknet_leaf_177_clk),
    .D(_01214_),
    .Q(\cur_mb_mem[132][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19917_ (.CLK(clknet_leaf_76_clk),
    .D(_01215_),
    .Q(\cur_mb_mem[133][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19918_ (.CLK(clknet_leaf_54_clk),
    .D(_01216_),
    .Q(\cur_mb_mem[133][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19919_ (.CLK(clknet_leaf_77_clk),
    .D(_01217_),
    .Q(\cur_mb_mem[133][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19920_ (.CLK(clknet_leaf_74_clk),
    .D(_01218_),
    .Q(\cur_mb_mem[133][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19921_ (.CLK(clknet_leaf_83_clk),
    .D(_01219_),
    .Q(\cur_mb_mem[133][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19922_ (.CLK(clknet_leaf_83_clk),
    .D(_01220_),
    .Q(\cur_mb_mem[133][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19923_ (.CLK(clknet_leaf_50_clk),
    .D(_01221_),
    .Q(\cur_mb_mem[133][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19924_ (.CLK(clknet_leaf_50_clk),
    .D(_01222_),
    .Q(\cur_mb_mem[133][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19925_ (.CLK(clknet_leaf_262_clk),
    .D(_01223_),
    .Q(\cur_mb_mem[134][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19926_ (.CLK(clknet_leaf_236_clk),
    .D(_01224_),
    .Q(\cur_mb_mem[134][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19927_ (.CLK(clknet_leaf_262_clk),
    .D(_01225_),
    .Q(\cur_mb_mem[134][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19928_ (.CLK(clknet_leaf_262_clk),
    .D(_01226_),
    .Q(\cur_mb_mem[134][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19929_ (.CLK(clknet_leaf_196_clk),
    .D(_01227_),
    .Q(\cur_mb_mem[134][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19930_ (.CLK(clknet_leaf_168_clk),
    .D(_01228_),
    .Q(\cur_mb_mem[134][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19931_ (.CLK(clknet_leaf_235_clk),
    .D(_01229_),
    .Q(\cur_mb_mem[134][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19932_ (.CLK(clknet_leaf_246_clk),
    .D(_01230_),
    .Q(\cur_mb_mem[134][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19933_ (.CLK(clknet_leaf_247_clk),
    .D(_01231_),
    .Q(\cur_mb_mem[135][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19934_ (.CLK(clknet_leaf_164_clk),
    .D(_01232_),
    .Q(\cur_mb_mem[135][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19935_ (.CLK(clknet_leaf_247_clk),
    .D(_01233_),
    .Q(\cur_mb_mem[135][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19936_ (.CLK(clknet_leaf_247_clk),
    .D(_01234_),
    .Q(\cur_mb_mem[135][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19937_ (.CLK(clknet_leaf_231_clk),
    .D(_01235_),
    .Q(\cur_mb_mem[135][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19938_ (.CLK(clknet_leaf_231_clk),
    .D(_01236_),
    .Q(\cur_mb_mem[135][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19939_ (.CLK(clknet_leaf_246_clk),
    .D(_01237_),
    .Q(\cur_mb_mem[135][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19940_ (.CLK(clknet_leaf_246_clk),
    .D(_01238_),
    .Q(\cur_mb_mem[135][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19941_ (.CLK(clknet_leaf_110_clk),
    .D(_01239_),
    .Q(\cur_mb_mem[136][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19942_ (.CLK(clknet_leaf_63_clk),
    .D(_01240_),
    .Q(\cur_mb_mem[136][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19943_ (.CLK(clknet_leaf_143_clk),
    .D(_01241_),
    .Q(\cur_mb_mem[136][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19944_ (.CLK(clknet_leaf_110_clk),
    .D(_01242_),
    .Q(\cur_mb_mem[136][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19945_ (.CLK(clknet_leaf_108_clk),
    .D(_01243_),
    .Q(\cur_mb_mem[136][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19946_ (.CLK(clknet_leaf_108_clk),
    .D(_01244_),
    .Q(\cur_mb_mem[136][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19947_ (.CLK(clknet_leaf_145_clk),
    .D(_01245_),
    .Q(\cur_mb_mem[136][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19948_ (.CLK(clknet_leaf_177_clk),
    .D(_01246_),
    .Q(\cur_mb_mem[136][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19949_ (.CLK(clknet_leaf_71_clk),
    .D(_01247_),
    .Q(\cur_mb_mem[137][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19950_ (.CLK(clknet_leaf_59_clk),
    .D(_01248_),
    .Q(\cur_mb_mem[137][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19951_ (.CLK(clknet_leaf_71_clk),
    .D(_01249_),
    .Q(\cur_mb_mem[137][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19952_ (.CLK(clknet_leaf_73_clk),
    .D(_01250_),
    .Q(\cur_mb_mem[137][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19953_ (.CLK(clknet_leaf_59_clk),
    .D(_01251_),
    .Q(\cur_mb_mem[137][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19954_ (.CLK(clknet_leaf_61_clk),
    .D(_01252_),
    .Q(\cur_mb_mem[137][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19955_ (.CLK(clknet_leaf_150_clk),
    .D(_01253_),
    .Q(\cur_mb_mem[137][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19956_ (.CLK(clknet_leaf_151_clk),
    .D(_01254_),
    .Q(\cur_mb_mem[137][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19957_ (.CLK(clknet_leaf_77_clk),
    .D(_01255_),
    .Q(\cur_mb_mem[138][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19958_ (.CLK(clknet_leaf_71_clk),
    .D(_01256_),
    .Q(\cur_mb_mem[138][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19959_ (.CLK(clknet_leaf_77_clk),
    .D(_01257_),
    .Q(\cur_mb_mem[138][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19960_ (.CLK(clknet_leaf_74_clk),
    .D(_01258_),
    .Q(\cur_mb_mem[138][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19961_ (.CLK(clknet_leaf_57_clk),
    .D(_01259_),
    .Q(\cur_mb_mem[138][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19962_ (.CLK(clknet_leaf_58_clk),
    .D(_01260_),
    .Q(\cur_mb_mem[138][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19963_ (.CLK(clknet_leaf_239_clk),
    .D(_01261_),
    .Q(\cur_mb_mem[138][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19964_ (.CLK(clknet_leaf_151_clk),
    .D(_01262_),
    .Q(\cur_mb_mem[138][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19965_ (.CLK(clknet_leaf_37_clk),
    .D(_01263_),
    .Q(\cur_mb_mem[139][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19966_ (.CLK(clknet_leaf_347_clk),
    .D(_01264_),
    .Q(\cur_mb_mem[139][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19967_ (.CLK(clknet_leaf_345_clk),
    .D(_01265_),
    .Q(\cur_mb_mem[139][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19968_ (.CLK(clknet_leaf_37_clk),
    .D(_01266_),
    .Q(\cur_mb_mem[139][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19969_ (.CLK(clknet_leaf_106_clk),
    .D(_01267_),
    .Q(\cur_mb_mem[139][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19970_ (.CLK(clknet_leaf_106_clk),
    .D(_01268_),
    .Q(\cur_mb_mem[139][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19971_ (.CLK(clknet_leaf_41_clk),
    .D(_01269_),
    .Q(\cur_mb_mem[139][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19972_ (.CLK(clknet_leaf_51_clk),
    .D(_01270_),
    .Q(\cur_mb_mem[139][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19973_ (.CLK(clknet_leaf_85_clk),
    .D(_01271_),
    .Q(\cur_mb_mem[140][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19974_ (.CLK(clknet_leaf_55_clk),
    .D(_01272_),
    .Q(\cur_mb_mem[140][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19975_ (.CLK(clknet_leaf_85_clk),
    .D(_01273_),
    .Q(\cur_mb_mem[140][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19976_ (.CLK(clknet_leaf_85_clk),
    .D(_01274_),
    .Q(\cur_mb_mem[140][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19977_ (.CLK(clknet_leaf_133_clk),
    .D(_01275_),
    .Q(\cur_mb_mem[140][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19978_ (.CLK(clknet_leaf_133_clk),
    .D(_01276_),
    .Q(\cur_mb_mem[140][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19979_ (.CLK(clknet_leaf_56_clk),
    .D(_01277_),
    .Q(\cur_mb_mem[140][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19980_ (.CLK(clknet_leaf_141_clk),
    .D(_01278_),
    .Q(\cur_mb_mem[140][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19981_ (.CLK(clknet_leaf_70_clk),
    .D(_01279_),
    .Q(\cur_mb_mem[141][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19982_ (.CLK(clknet_leaf_55_clk),
    .D(_01280_),
    .Q(\cur_mb_mem[141][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19983_ (.CLK(clknet_leaf_46_clk),
    .D(_01281_),
    .Q(\cur_mb_mem[141][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19984_ (.CLK(clknet_leaf_30_clk),
    .D(_01282_),
    .Q(\cur_mb_mem[141][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19985_ (.CLK(clknet_leaf_134_clk),
    .D(_01283_),
    .Q(\cur_mb_mem[141][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19986_ (.CLK(clknet_leaf_134_clk),
    .D(_01284_),
    .Q(\cur_mb_mem[141][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19987_ (.CLK(clknet_leaf_41_clk),
    .D(_01285_),
    .Q(\cur_mb_mem[141][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19988_ (.CLK(clknet_leaf_42_clk),
    .D(_01286_),
    .Q(\cur_mb_mem[141][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19989_ (.CLK(clknet_leaf_347_clk),
    .D(_01287_),
    .Q(\cur_mb_mem[142][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19990_ (.CLK(clknet_leaf_347_clk),
    .D(_01288_),
    .Q(\cur_mb_mem[142][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19991_ (.CLK(clknet_leaf_345_clk),
    .D(_01289_),
    .Q(\cur_mb_mem[142][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19992_ (.CLK(clknet_leaf_38_clk),
    .D(_01290_),
    .Q(\cur_mb_mem[142][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19993_ (.CLK(clknet_leaf_38_clk),
    .D(_01291_),
    .Q(\cur_mb_mem[142][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19994_ (.CLK(clknet_leaf_38_clk),
    .D(_01292_),
    .Q(\cur_mb_mem[142][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19995_ (.CLK(clknet_leaf_46_clk),
    .D(_01293_),
    .Q(\cur_mb_mem[142][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19996_ (.CLK(clknet_leaf_61_clk),
    .D(_01294_),
    .Q(\cur_mb_mem[142][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19997_ (.CLK(clknet_leaf_260_clk),
    .D(_01295_),
    .Q(\cur_mb_mem[143][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19998_ (.CLK(clknet_leaf_327_clk),
    .D(_01296_),
    .Q(\cur_mb_mem[143][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19999_ (.CLK(clknet_leaf_260_clk),
    .D(_01297_),
    .Q(\cur_mb_mem[143][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20000_ (.CLK(clknet_leaf_260_clk),
    .D(_01298_),
    .Q(\cur_mb_mem[143][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20001_ (.CLK(clknet_leaf_28_clk),
    .D(_01299_),
    .Q(\cur_mb_mem[143][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20002_ (.CLK(clknet_leaf_27_clk),
    .D(_01300_),
    .Q(\cur_mb_mem[143][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20003_ (.CLK(clknet_leaf_70_clk),
    .D(_01301_),
    .Q(\cur_mb_mem[143][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20004_ (.CLK(clknet_leaf_237_clk),
    .D(_01302_),
    .Q(\cur_mb_mem[143][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20005_ (.CLK(clknet_leaf_260_clk),
    .D(_01303_),
    .Q(\cur_mb_mem[144][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20006_ (.CLK(clknet_leaf_39_clk),
    .D(_01304_),
    .Q(\cur_mb_mem[144][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20007_ (.CLK(clknet_leaf_260_clk),
    .D(_01305_),
    .Q(\cur_mb_mem[144][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20008_ (.CLK(clknet_leaf_260_clk),
    .D(_01306_),
    .Q(\cur_mb_mem[144][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20009_ (.CLK(clknet_leaf_11_clk),
    .D(_01307_),
    .Q(\cur_mb_mem[144][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20010_ (.CLK(clknet_leaf_11_clk),
    .D(_01308_),
    .Q(\cur_mb_mem[144][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20011_ (.CLK(clknet_leaf_329_clk),
    .D(_01309_),
    .Q(\cur_mb_mem[144][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20012_ (.CLK(clknet_leaf_41_clk),
    .D(_01310_),
    .Q(\cur_mb_mem[144][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20013_ (.CLK(clknet_leaf_8_clk),
    .D(_01311_),
    .Q(\cur_mb_mem[145][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20014_ (.CLK(clknet_leaf_346_clk),
    .D(_01312_),
    .Q(\cur_mb_mem[145][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20015_ (.CLK(clknet_leaf_346_clk),
    .D(_01313_),
    .Q(\cur_mb_mem[145][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20016_ (.CLK(clknet_leaf_7_clk),
    .D(_01314_),
    .Q(\cur_mb_mem[145][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20017_ (.CLK(clknet_leaf_25_clk),
    .D(_01315_),
    .Q(\cur_mb_mem[145][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20018_ (.CLK(clknet_leaf_25_clk),
    .D(_01316_),
    .Q(\cur_mb_mem[145][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20019_ (.CLK(clknet_leaf_42_clk),
    .D(_01317_),
    .Q(\cur_mb_mem[145][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20020_ (.CLK(clknet_leaf_42_clk),
    .D(_01318_),
    .Q(\cur_mb_mem[145][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20021_ (.CLK(clknet_leaf_32_clk),
    .D(_01319_),
    .Q(\cur_mb_mem[146][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20022_ (.CLK(clknet_leaf_35_clk),
    .D(_01320_),
    .Q(\cur_mb_mem[146][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20023_ (.CLK(clknet_leaf_41_clk),
    .D(_01321_),
    .Q(\cur_mb_mem[146][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20024_ (.CLK(clknet_leaf_20_clk),
    .D(_01322_),
    .Q(\cur_mb_mem[146][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20025_ (.CLK(clknet_leaf_78_clk),
    .D(_01323_),
    .Q(\cur_mb_mem[146][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20026_ (.CLK(clknet_leaf_78_clk),
    .D(_01324_),
    .Q(\cur_mb_mem[146][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20027_ (.CLK(clknet_leaf_29_clk),
    .D(_01325_),
    .Q(\cur_mb_mem[146][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20028_ (.CLK(clknet_leaf_56_clk),
    .D(_01326_),
    .Q(\cur_mb_mem[146][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20029_ (.CLK(clknet_leaf_90_clk),
    .D(_01327_),
    .Q(\cur_mb_mem[147][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20030_ (.CLK(clknet_leaf_36_clk),
    .D(_01328_),
    .Q(\cur_mb_mem[147][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20031_ (.CLK(clknet_leaf_87_clk),
    .D(_01329_),
    .Q(\cur_mb_mem[147][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20032_ (.CLK(clknet_leaf_77_clk),
    .D(_01330_),
    .Q(\cur_mb_mem[147][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20033_ (.CLK(clknet_leaf_16_clk),
    .D(_01331_),
    .Q(\cur_mb_mem[147][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20034_ (.CLK(clknet_leaf_16_clk),
    .D(_01332_),
    .Q(\cur_mb_mem[147][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20035_ (.CLK(clknet_leaf_333_clk),
    .D(_01333_),
    .Q(\cur_mb_mem[147][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20036_ (.CLK(clknet_leaf_328_clk),
    .D(_01334_),
    .Q(\cur_mb_mem[147][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20037_ (.CLK(clknet_leaf_88_clk),
    .D(_01335_),
    .Q(\cur_mb_mem[148][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20038_ (.CLK(clknet_leaf_31_clk),
    .D(_01336_),
    .Q(\cur_mb_mem[148][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20039_ (.CLK(clknet_leaf_88_clk),
    .D(_01337_),
    .Q(\cur_mb_mem[148][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20040_ (.CLK(clknet_leaf_88_clk),
    .D(_01338_),
    .Q(\cur_mb_mem[148][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20041_ (.CLK(clknet_leaf_58_clk),
    .D(_01339_),
    .Q(\cur_mb_mem[148][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20042_ (.CLK(clknet_leaf_57_clk),
    .D(_01340_),
    .Q(\cur_mb_mem[148][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20043_ (.CLK(clknet_leaf_56_clk),
    .D(_01341_),
    .Q(\cur_mb_mem[148][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20044_ (.CLK(clknet_leaf_61_clk),
    .D(_01342_),
    .Q(\cur_mb_mem[148][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20045_ (.CLK(clknet_leaf_0_clk),
    .D(_01343_),
    .Q(\cur_mb_mem[149][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20046_ (.CLK(clknet_leaf_26_clk),
    .D(_01344_),
    .Q(\cur_mb_mem[149][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20047_ (.CLK(clknet_leaf_0_clk),
    .D(_01345_),
    .Q(\cur_mb_mem[149][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20048_ (.CLK(clknet_leaf_2_clk),
    .D(_01346_),
    .Q(\cur_mb_mem[149][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20049_ (.CLK(clknet_leaf_12_clk),
    .D(_01347_),
    .Q(\cur_mb_mem[149][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20050_ (.CLK(clknet_leaf_12_clk),
    .D(_01348_),
    .Q(\cur_mb_mem[149][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20051_ (.CLK(clknet_leaf_19_clk),
    .D(_01349_),
    .Q(\cur_mb_mem[149][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20052_ (.CLK(clknet_leaf_34_clk),
    .D(_01350_),
    .Q(\cur_mb_mem[149][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20053_ (.CLK(clknet_leaf_6_clk),
    .D(_01351_),
    .Q(\cur_mb_mem[150][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20054_ (.CLK(clknet_leaf_39_clk),
    .D(_01352_),
    .Q(\cur_mb_mem[150][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20055_ (.CLK(clknet_leaf_6_clk),
    .D(_01353_),
    .Q(\cur_mb_mem[150][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20056_ (.CLK(clknet_leaf_381_clk),
    .D(_01354_),
    .Q(\cur_mb_mem[150][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20057_ (.CLK(clknet_leaf_13_clk),
    .D(_01355_),
    .Q(\cur_mb_mem[150][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20058_ (.CLK(clknet_leaf_0_clk),
    .D(_01356_),
    .Q(\cur_mb_mem[150][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20059_ (.CLK(clknet_leaf_326_clk),
    .D(_01357_),
    .Q(\cur_mb_mem[150][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20060_ (.CLK(clknet_leaf_322_clk),
    .D(_01358_),
    .Q(\cur_mb_mem[150][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20061_ (.CLK(clknet_leaf_9_clk),
    .D(_01359_),
    .Q(\cur_mb_mem[151][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20062_ (.CLK(clknet_leaf_345_clk),
    .D(_01360_),
    .Q(\cur_mb_mem[151][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20063_ (.CLK(clknet_leaf_12_clk),
    .D(_01361_),
    .Q(\cur_mb_mem[151][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20064_ (.CLK(clknet_leaf_9_clk),
    .D(_01362_),
    .Q(\cur_mb_mem[151][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20065_ (.CLK(clknet_leaf_14_clk),
    .D(_01363_),
    .Q(\cur_mb_mem[151][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20066_ (.CLK(clknet_leaf_15_clk),
    .D(_01364_),
    .Q(\cur_mb_mem[151][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20067_ (.CLK(clknet_leaf_326_clk),
    .D(_01365_),
    .Q(\cur_mb_mem[151][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20068_ (.CLK(clknet_leaf_322_clk),
    .D(_01366_),
    .Q(\cur_mb_mem[151][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20069_ (.CLK(clknet_leaf_72_clk),
    .D(_01367_),
    .Q(\cur_mb_mem[152][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20070_ (.CLK(clknet_leaf_57_clk),
    .D(_01368_),
    .Q(\cur_mb_mem[152][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20071_ (.CLK(clknet_leaf_72_clk),
    .D(_01369_),
    .Q(\cur_mb_mem[152][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20072_ (.CLK(clknet_leaf_73_clk),
    .D(_01370_),
    .Q(\cur_mb_mem[152][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20073_ (.CLK(clknet_leaf_24_clk),
    .D(_01371_),
    .Q(\cur_mb_mem[152][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20074_ (.CLK(clknet_leaf_24_clk),
    .D(_01372_),
    .Q(\cur_mb_mem[152][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20075_ (.CLK(clknet_leaf_48_clk),
    .D(_01373_),
    .Q(\cur_mb_mem[152][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20076_ (.CLK(clknet_leaf_48_clk),
    .D(_01374_),
    .Q(\cur_mb_mem[152][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20077_ (.CLK(clknet_leaf_90_clk),
    .D(_01375_),
    .Q(\cur_mb_mem[153][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20078_ (.CLK(clknet_leaf_19_clk),
    .D(_01376_),
    .Q(\cur_mb_mem[153][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20079_ (.CLK(clknet_leaf_90_clk),
    .D(_01377_),
    .Q(\cur_mb_mem[153][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20080_ (.CLK(clknet_leaf_26_clk),
    .D(_01378_),
    .Q(\cur_mb_mem[153][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20081_ (.CLK(clknet_leaf_25_clk),
    .D(_01379_),
    .Q(\cur_mb_mem[153][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20082_ (.CLK(clknet_leaf_25_clk),
    .D(_01380_),
    .Q(\cur_mb_mem[153][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20083_ (.CLK(clknet_leaf_10_clk),
    .D(_01381_),
    .Q(\cur_mb_mem[153][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20084_ (.CLK(clknet_leaf_27_clk),
    .D(_01382_),
    .Q(\cur_mb_mem[153][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20085_ (.CLK(clknet_leaf_3_clk),
    .D(_01383_),
    .Q(\cur_mb_mem[154][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20086_ (.CLK(clknet_leaf_26_clk),
    .D(_01384_),
    .Q(\cur_mb_mem[154][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20087_ (.CLK(clknet_leaf_2_clk),
    .D(_01385_),
    .Q(\cur_mb_mem[154][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20088_ (.CLK(clknet_leaf_3_clk),
    .D(_01386_),
    .Q(\cur_mb_mem[154][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20089_ (.CLK(clknet_leaf_24_clk),
    .D(_01387_),
    .Q(\cur_mb_mem[154][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20090_ (.CLK(clknet_leaf_25_clk),
    .D(_01388_),
    .Q(\cur_mb_mem[154][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20091_ (.CLK(clknet_leaf_18_clk),
    .D(_01389_),
    .Q(\cur_mb_mem[154][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20092_ (.CLK(clknet_leaf_27_clk),
    .D(_01390_),
    .Q(\cur_mb_mem[154][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20093_ (.CLK(clknet_leaf_31_clk),
    .D(_01391_),
    .Q(\cur_mb_mem[155][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20094_ (.CLK(clknet_leaf_43_clk),
    .D(_01392_),
    .Q(\cur_mb_mem[155][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20095_ (.CLK(clknet_leaf_24_clk),
    .D(_01393_),
    .Q(\cur_mb_mem[155][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20096_ (.CLK(clknet_leaf_31_clk),
    .D(_01394_),
    .Q(\cur_mb_mem[155][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20097_ (.CLK(clknet_leaf_20_clk),
    .D(_01395_),
    .Q(\cur_mb_mem[155][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20098_ (.CLK(clknet_leaf_22_clk),
    .D(_01396_),
    .Q(\cur_mb_mem[155][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20099_ (.CLK(clknet_leaf_43_clk),
    .D(_01397_),
    .Q(\cur_mb_mem[155][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20100_ (.CLK(clknet_leaf_43_clk),
    .D(_01398_),
    .Q(\cur_mb_mem[155][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20101_ (.CLK(clknet_leaf_0_clk),
    .D(_01399_),
    .Q(\cur_mb_mem[156][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20102_ (.CLK(clknet_leaf_26_clk),
    .D(_01400_),
    .Q(\cur_mb_mem[156][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20103_ (.CLK(clknet_leaf_0_clk),
    .D(_01401_),
    .Q(\cur_mb_mem[156][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20104_ (.CLK(clknet_leaf_0_clk),
    .D(_01402_),
    .Q(\cur_mb_mem[156][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20105_ (.CLK(clknet_leaf_14_clk),
    .D(_01403_),
    .Q(\cur_mb_mem[156][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20106_ (.CLK(clknet_leaf_0_clk),
    .D(_01404_),
    .Q(\cur_mb_mem[156][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20107_ (.CLK(clknet_leaf_20_clk),
    .D(_01405_),
    .Q(\cur_mb_mem[156][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20108_ (.CLK(clknet_leaf_34_clk),
    .D(_01406_),
    .Q(\cur_mb_mem[156][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20109_ (.CLK(clknet_leaf_2_clk),
    .D(_01407_),
    .Q(\cur_mb_mem[157][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20110_ (.CLK(clknet_leaf_36_clk),
    .D(_01408_),
    .Q(\cur_mb_mem[157][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20111_ (.CLK(clknet_leaf_1_clk),
    .D(_01409_),
    .Q(\cur_mb_mem[157][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20112_ (.CLK(clknet_leaf_2_clk),
    .D(_01410_),
    .Q(\cur_mb_mem[157][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20113_ (.CLK(clknet_leaf_26_clk),
    .D(_01411_),
    .Q(\cur_mb_mem[157][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20114_ (.CLK(clknet_leaf_26_clk),
    .D(_01412_),
    .Q(\cur_mb_mem[157][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20115_ (.CLK(clknet_leaf_326_clk),
    .D(_01413_),
    .Q(\cur_mb_mem[157][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20116_ (.CLK(clknet_leaf_328_clk),
    .D(_01414_),
    .Q(\cur_mb_mem[157][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20117_ (.CLK(clknet_leaf_13_clk),
    .D(_01415_),
    .Q(\cur_mb_mem[158][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20118_ (.CLK(clknet_leaf_38_clk),
    .D(_01416_),
    .Q(\cur_mb_mem[158][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20119_ (.CLK(clknet_leaf_19_clk),
    .D(_01417_),
    .Q(\cur_mb_mem[158][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20120_ (.CLK(clknet_leaf_7_clk),
    .D(_01418_),
    .Q(\cur_mb_mem[158][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20121_ (.CLK(clknet_leaf_15_clk),
    .D(_01419_),
    .Q(\cur_mb_mem[158][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20122_ (.CLK(clknet_leaf_15_clk),
    .D(_01420_),
    .Q(\cur_mb_mem[158][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20123_ (.CLK(clknet_leaf_39_clk),
    .D(_01421_),
    .Q(\cur_mb_mem[158][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20124_ (.CLK(clknet_leaf_39_clk),
    .D(_01422_),
    .Q(\cur_mb_mem[158][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20125_ (.CLK(clknet_leaf_165_clk),
    .D(_01423_),
    .Q(\cur_mb_mem[159][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20126_ (.CLK(clknet_leaf_240_clk),
    .D(_01424_),
    .Q(\cur_mb_mem[159][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20127_ (.CLK(clknet_leaf_165_clk),
    .D(_01425_),
    .Q(\cur_mb_mem[159][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20128_ (.CLK(clknet_leaf_165_clk),
    .D(_01426_),
    .Q(\cur_mb_mem[159][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20129_ (.CLK(clknet_leaf_25_clk),
    .D(_01427_),
    .Q(\cur_mb_mem[159][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20130_ (.CLK(clknet_leaf_77_clk),
    .D(_01428_),
    .Q(\cur_mb_mem[159][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20131_ (.CLK(clknet_leaf_163_clk),
    .D(_01429_),
    .Q(\cur_mb_mem[159][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20132_ (.CLK(clknet_leaf_243_clk),
    .D(_01430_),
    .Q(\cur_mb_mem[159][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20133_ (.CLK(clknet_leaf_174_clk),
    .D(_01431_),
    .Q(\cur_mb_mem[160][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20134_ (.CLK(clknet_leaf_337_clk),
    .D(_01432_),
    .Q(\cur_mb_mem[160][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20135_ (.CLK(clknet_leaf_166_clk),
    .D(_01433_),
    .Q(\cur_mb_mem[160][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20136_ (.CLK(clknet_leaf_166_clk),
    .D(_01434_),
    .Q(\cur_mb_mem[160][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20137_ (.CLK(clknet_leaf_45_clk),
    .D(_01435_),
    .Q(\cur_mb_mem[160][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20138_ (.CLK(clknet_leaf_45_clk),
    .D(_01436_),
    .Q(\cur_mb_mem[160][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20139_ (.CLK(clknet_leaf_232_clk),
    .D(_01437_),
    .Q(\cur_mb_mem[160][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20140_ (.CLK(clknet_leaf_163_clk),
    .D(_01438_),
    .Q(\cur_mb_mem[160][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20141_ (.CLK(clknet_leaf_147_clk),
    .D(_01439_),
    .Q(\cur_mb_mem[161][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20142_ (.CLK(clknet_leaf_326_clk),
    .D(_01440_),
    .Q(\cur_mb_mem[161][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20143_ (.CLK(clknet_leaf_157_clk),
    .D(_01441_),
    .Q(\cur_mb_mem[161][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20144_ (.CLK(clknet_leaf_140_clk),
    .D(_01442_),
    .Q(\cur_mb_mem[161][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20145_ (.CLK(clknet_leaf_60_clk),
    .D(_01443_),
    .Q(\cur_mb_mem[161][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20146_ (.CLK(clknet_leaf_55_clk),
    .D(_01444_),
    .Q(\cur_mb_mem[161][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20147_ (.CLK(clknet_leaf_334_clk),
    .D(_01445_),
    .Q(\cur_mb_mem[161][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20148_ (.CLK(clknet_leaf_241_clk),
    .D(_01446_),
    .Q(\cur_mb_mem[161][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20149_ (.CLK(clknet_leaf_316_clk),
    .D(_01447_),
    .Q(\cur_mb_mem[162][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20150_ (.CLK(clknet_leaf_329_clk),
    .D(_01448_),
    .Q(\cur_mb_mem[162][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20151_ (.CLK(clknet_leaf_315_clk),
    .D(_01449_),
    .Q(\cur_mb_mem[162][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20152_ (.CLK(clknet_leaf_254_clk),
    .D(_01450_),
    .Q(\cur_mb_mem[162][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20153_ (.CLK(clknet_leaf_331_clk),
    .D(_01451_),
    .Q(\cur_mb_mem[162][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20154_ (.CLK(clknet_leaf_331_clk),
    .D(_01452_),
    .Q(\cur_mb_mem[162][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20155_ (.CLK(clknet_leaf_146_clk),
    .D(_01453_),
    .Q(\cur_mb_mem[162][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20156_ (.CLK(clknet_leaf_146_clk),
    .D(_01454_),
    .Q(\cur_mb_mem[162][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20157_ (.CLK(clknet_leaf_88_clk),
    .D(_01455_),
    .Q(\cur_mb_mem[163][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20158_ (.CLK(clknet_leaf_62_clk),
    .D(_01456_),
    .Q(\cur_mb_mem[163][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20159_ (.CLK(clknet_leaf_88_clk),
    .D(_01457_),
    .Q(\cur_mb_mem[163][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20160_ (.CLK(clknet_leaf_93_clk),
    .D(_01458_),
    .Q(\cur_mb_mem[163][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20161_ (.CLK(clknet_leaf_60_clk),
    .D(_01459_),
    .Q(\cur_mb_mem[163][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20162_ (.CLK(clknet_leaf_56_clk),
    .D(_01460_),
    .Q(\cur_mb_mem[163][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20163_ (.CLK(clknet_leaf_244_clk),
    .D(_01461_),
    .Q(\cur_mb_mem[163][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20164_ (.CLK(clknet_leaf_239_clk),
    .D(_01462_),
    .Q(\cur_mb_mem[163][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20165_ (.CLK(clknet_leaf_263_clk),
    .D(_01463_),
    .Q(\cur_mb_mem[164][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20166_ (.CLK(clknet_leaf_336_clk),
    .D(_01464_),
    .Q(\cur_mb_mem[164][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20167_ (.CLK(clknet_leaf_263_clk),
    .D(_01465_),
    .Q(\cur_mb_mem[164][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20168_ (.CLK(clknet_leaf_263_clk),
    .D(_01466_),
    .Q(\cur_mb_mem[164][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20169_ (.CLK(clknet_leaf_178_clk),
    .D(_01467_),
    .Q(\cur_mb_mem[164][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20170_ (.CLK(clknet_leaf_178_clk),
    .D(_01468_),
    .Q(\cur_mb_mem[164][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20171_ (.CLK(clknet_leaf_332_clk),
    .D(_01469_),
    .Q(\cur_mb_mem[164][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20172_ (.CLK(clknet_leaf_175_clk),
    .D(_01470_),
    .Q(\cur_mb_mem[164][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20173_ (.CLK(clknet_leaf_84_clk),
    .D(_01471_),
    .Q(\cur_mb_mem[165][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20174_ (.CLK(clknet_leaf_62_clk),
    .D(_01472_),
    .Q(\cur_mb_mem[165][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20175_ (.CLK(clknet_leaf_90_clk),
    .D(_01473_),
    .Q(\cur_mb_mem[165][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20176_ (.CLK(clknet_leaf_91_clk),
    .D(_01474_),
    .Q(\cur_mb_mem[165][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20177_ (.CLK(clknet_leaf_44_clk),
    .D(_01475_),
    .Q(\cur_mb_mem[165][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20178_ (.CLK(clknet_leaf_45_clk),
    .D(_01476_),
    .Q(\cur_mb_mem[165][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20179_ (.CLK(clknet_leaf_158_clk),
    .D(_01477_),
    .Q(\cur_mb_mem[165][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20180_ (.CLK(clknet_leaf_333_clk),
    .D(_01478_),
    .Q(\cur_mb_mem[165][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20181_ (.CLK(clknet_leaf_161_clk),
    .D(_01479_),
    .Q(\cur_mb_mem[166][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20182_ (.CLK(clknet_leaf_348_clk),
    .D(_01480_),
    .Q(\cur_mb_mem[166][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20183_ (.CLK(clknet_leaf_161_clk),
    .D(_01481_),
    .Q(\cur_mb_mem[166][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20184_ (.CLK(clknet_leaf_175_clk),
    .D(_01482_),
    .Q(\cur_mb_mem[166][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20185_ (.CLK(clknet_leaf_377_clk),
    .D(_01483_),
    .Q(\cur_mb_mem[166][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20186_ (.CLK(clknet_leaf_377_clk),
    .D(_01484_),
    .Q(\cur_mb_mem[166][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20187_ (.CLK(clknet_leaf_349_clk),
    .D(_01485_),
    .Q(\cur_mb_mem[166][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20188_ (.CLK(clknet_leaf_242_clk),
    .D(_01486_),
    .Q(\cur_mb_mem[166][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20189_ (.CLK(clknet_leaf_252_clk),
    .D(_01487_),
    .Q(\cur_mb_mem[167][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20190_ (.CLK(clknet_leaf_316_clk),
    .D(_01488_),
    .Q(\cur_mb_mem[167][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20191_ (.CLK(clknet_leaf_252_clk),
    .D(_01489_),
    .Q(\cur_mb_mem[167][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20192_ (.CLK(clknet_leaf_318_clk),
    .D(_01490_),
    .Q(\cur_mb_mem[167][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20193_ (.CLK(clknet_leaf_332_clk),
    .D(_01491_),
    .Q(\cur_mb_mem[167][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20194_ (.CLK(clknet_leaf_329_clk),
    .D(_01492_),
    .Q(\cur_mb_mem[167][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20195_ (.CLK(clknet_leaf_327_clk),
    .D(_01493_),
    .Q(\cur_mb_mem[167][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20196_ (.CLK(clknet_leaf_320_clk),
    .D(_01494_),
    .Q(\cur_mb_mem[167][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20197_ (.CLK(clknet_leaf_70_clk),
    .D(_01495_),
    .Q(\cur_mb_mem[168][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20198_ (.CLK(clknet_leaf_335_clk),
    .D(_01496_),
    .Q(\cur_mb_mem[168][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20199_ (.CLK(clknet_leaf_69_clk),
    .D(_01497_),
    .Q(\cur_mb_mem[168][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20200_ (.CLK(clknet_leaf_67_clk),
    .D(_01498_),
    .Q(\cur_mb_mem[168][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20201_ (.CLK(clknet_leaf_51_clk),
    .D(_01499_),
    .Q(\cur_mb_mem[168][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20202_ (.CLK(clknet_leaf_40_clk),
    .D(_01500_),
    .Q(\cur_mb_mem[168][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20203_ (.CLK(clknet_leaf_147_clk),
    .D(_01501_),
    .Q(\cur_mb_mem[168][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20204_ (.CLK(clknet_leaf_48_clk),
    .D(_01502_),
    .Q(\cur_mb_mem[168][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20205_ (.CLK(clknet_leaf_70_clk),
    .D(_01503_),
    .Q(\cur_mb_mem[169][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20206_ (.CLK(clknet_leaf_57_clk),
    .D(_01504_),
    .Q(\cur_mb_mem[169][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20207_ (.CLK(clknet_leaf_68_clk),
    .D(_01505_),
    .Q(\cur_mb_mem[169][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20208_ (.CLK(clknet_leaf_67_clk),
    .D(_01506_),
    .Q(\cur_mb_mem[169][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20209_ (.CLK(clknet_leaf_381_clk),
    .D(_01507_),
    .Q(\cur_mb_mem[169][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20210_ (.CLK(clknet_leaf_379_clk),
    .D(_01508_),
    .Q(\cur_mb_mem[169][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20211_ (.CLK(clknet_leaf_60_clk),
    .D(_01509_),
    .Q(\cur_mb_mem[169][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20212_ (.CLK(clknet_leaf_345_clk),
    .D(_01510_),
    .Q(\cur_mb_mem[169][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20213_ (.CLK(clknet_leaf_65_clk),
    .D(_01511_),
    .Q(\cur_mb_mem[170][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20214_ (.CLK(clknet_leaf_56_clk),
    .D(_01512_),
    .Q(\cur_mb_mem[170][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20215_ (.CLK(clknet_leaf_142_clk),
    .D(_01513_),
    .Q(\cur_mb_mem[170][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20216_ (.CLK(clknet_leaf_65_clk),
    .D(_01514_),
    .Q(\cur_mb_mem[170][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20217_ (.CLK(clknet_leaf_377_clk),
    .D(_01515_),
    .Q(\cur_mb_mem[170][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20218_ (.CLK(clknet_leaf_350_clk),
    .D(_01516_),
    .Q(\cur_mb_mem[170][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20219_ (.CLK(clknet_leaf_339_clk),
    .D(_01517_),
    .Q(\cur_mb_mem[170][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20220_ (.CLK(clknet_leaf_335_clk),
    .D(_01518_),
    .Q(\cur_mb_mem[170][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20221_ (.CLK(clknet_leaf_67_clk),
    .D(_01519_),
    .Q(\cur_mb_mem[171][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20222_ (.CLK(clknet_leaf_354_clk),
    .D(_01520_),
    .Q(\cur_mb_mem[171][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20223_ (.CLK(clknet_leaf_67_clk),
    .D(_01521_),
    .Q(\cur_mb_mem[171][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20224_ (.CLK(clknet_leaf_66_clk),
    .D(_01522_),
    .Q(\cur_mb_mem[171][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20225_ (.CLK(clknet_leaf_349_clk),
    .D(_01523_),
    .Q(\cur_mb_mem[171][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20226_ (.CLK(clknet_leaf_349_clk),
    .D(_01524_),
    .Q(\cur_mb_mem[171][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20227_ (.CLK(clknet_leaf_352_clk),
    .D(_01525_),
    .Q(\cur_mb_mem[171][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20228_ (.CLK(clknet_leaf_152_clk),
    .D(_01526_),
    .Q(\cur_mb_mem[171][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20229_ (.CLK(clknet_leaf_67_clk),
    .D(_01527_),
    .Q(\cur_mb_mem[172][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20230_ (.CLK(clknet_leaf_324_clk),
    .D(_01528_),
    .Q(\cur_mb_mem[172][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20231_ (.CLK(clknet_leaf_94_clk),
    .D(_01529_),
    .Q(\cur_mb_mem[172][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20232_ (.CLK(clknet_leaf_92_clk),
    .D(_01530_),
    .Q(\cur_mb_mem[172][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20233_ (.CLK(clknet_leaf_357_clk),
    .D(_01531_),
    .Q(\cur_mb_mem[172][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20234_ (.CLK(clknet_leaf_305_clk),
    .D(_01532_),
    .Q(\cur_mb_mem[172][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20235_ (.CLK(clknet_leaf_157_clk),
    .D(_01533_),
    .Q(\cur_mb_mem[172][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20236_ (.CLK(clknet_leaf_152_clk),
    .D(_01534_),
    .Q(\cur_mb_mem[172][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20237_ (.CLK(clknet_leaf_37_clk),
    .D(_01535_),
    .Q(\cur_mb_mem[173][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20238_ (.CLK(clknet_leaf_38_clk),
    .D(_01536_),
    .Q(\cur_mb_mem[173][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20239_ (.CLK(clknet_leaf_348_clk),
    .D(_01537_),
    .Q(\cur_mb_mem[173][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20240_ (.CLK(clknet_leaf_38_clk),
    .D(_01538_),
    .Q(\cur_mb_mem[173][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20241_ (.CLK(clknet_leaf_352_clk),
    .D(_01539_),
    .Q(\cur_mb_mem[173][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20242_ (.CLK(clknet_leaf_379_clk),
    .D(_01540_),
    .Q(\cur_mb_mem[173][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20243_ (.CLK(clknet_leaf_47_clk),
    .D(_01541_),
    .Q(\cur_mb_mem[173][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20244_ (.CLK(clknet_leaf_343_clk),
    .D(_01542_),
    .Q(\cur_mb_mem[173][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20245_ (.CLK(clknet_leaf_381_clk),
    .D(_01543_),
    .Q(\cur_mb_mem[174][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20246_ (.CLK(clknet_leaf_338_clk),
    .D(_01544_),
    .Q(\cur_mb_mem[174][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20247_ (.CLK(clknet_leaf_380_clk),
    .D(_01545_),
    .Q(\cur_mb_mem[174][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20248_ (.CLK(clknet_leaf_381_clk),
    .D(_01546_),
    .Q(\cur_mb_mem[174][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20249_ (.CLK(clknet_leaf_356_clk),
    .D(_01547_),
    .Q(\cur_mb_mem[174][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20250_ (.CLK(clknet_leaf_350_clk),
    .D(_01548_),
    .Q(\cur_mb_mem[174][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20251_ (.CLK(clknet_leaf_332_clk),
    .D(_01549_),
    .Q(\cur_mb_mem[174][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20252_ (.CLK(clknet_leaf_332_clk),
    .D(_01550_),
    .Q(\cur_mb_mem[174][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20253_ (.CLK(clknet_leaf_311_clk),
    .D(_01551_),
    .Q(\cur_mb_mem[175][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20254_ (.CLK(clknet_leaf_355_clk),
    .D(_01552_),
    .Q(\cur_mb_mem[175][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20255_ (.CLK(clknet_leaf_312_clk),
    .D(_01553_),
    .Q(\cur_mb_mem[175][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20256_ (.CLK(clknet_leaf_311_clk),
    .D(_01554_),
    .Q(\cur_mb_mem[175][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20257_ (.CLK(clknet_leaf_55_clk),
    .D(_01555_),
    .Q(\cur_mb_mem[175][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20258_ (.CLK(clknet_leaf_55_clk),
    .D(_01556_),
    .Q(\cur_mb_mem[175][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20259_ (.CLK(clknet_leaf_151_clk),
    .D(_01557_),
    .Q(\cur_mb_mem[175][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20260_ (.CLK(clknet_leaf_334_clk),
    .D(_01558_),
    .Q(\cur_mb_mem[175][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20261_ (.CLK(clknet_leaf_168_clk),
    .D(_01559_),
    .Q(\cur_mb_mem[176][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20262_ (.CLK(clknet_leaf_155_clk),
    .D(_01560_),
    .Q(\cur_mb_mem[176][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20263_ (.CLK(clknet_leaf_167_clk),
    .D(_01561_),
    .Q(\cur_mb_mem[176][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20264_ (.CLK(clknet_leaf_168_clk),
    .D(_01562_),
    .Q(\cur_mb_mem[176][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20265_ (.CLK(clknet_leaf_192_clk),
    .D(_01563_),
    .Q(\cur_mb_mem[176][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20266_ (.CLK(clknet_leaf_172_clk),
    .D(_01564_),
    .Q(\cur_mb_mem[176][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20267_ (.CLK(clknet_leaf_160_clk),
    .D(_01565_),
    .Q(\cur_mb_mem[176][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20268_ (.CLK(clknet_leaf_153_clk),
    .D(_01566_),
    .Q(\cur_mb_mem[176][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20269_ (.CLK(clknet_leaf_272_clk),
    .D(_01567_),
    .Q(\cur_mb_mem[177][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20270_ (.CLK(clknet_leaf_236_clk),
    .D(_01568_),
    .Q(\cur_mb_mem[177][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20271_ (.CLK(clknet_leaf_272_clk),
    .D(_01569_),
    .Q(\cur_mb_mem[177][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20272_ (.CLK(clknet_leaf_270_clk),
    .D(_01570_),
    .Q(\cur_mb_mem[177][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20273_ (.CLK(clknet_leaf_230_clk),
    .D(_01571_),
    .Q(\cur_mb_mem[177][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20274_ (.CLK(clknet_leaf_230_clk),
    .D(_01572_),
    .Q(\cur_mb_mem[177][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20275_ (.CLK(clknet_leaf_244_clk),
    .D(_01573_),
    .Q(\cur_mb_mem[177][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20276_ (.CLK(clknet_leaf_156_clk),
    .D(_01574_),
    .Q(\cur_mb_mem[177][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20277_ (.CLK(clknet_leaf_63_clk),
    .D(_01575_),
    .Q(\cur_mb_mem[178][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20278_ (.CLK(clknet_leaf_63_clk),
    .D(_01576_),
    .Q(\cur_mb_mem[178][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20279_ (.CLK(clknet_leaf_63_clk),
    .D(_01577_),
    .Q(\cur_mb_mem[178][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20280_ (.CLK(clknet_leaf_66_clk),
    .D(_01578_),
    .Q(\cur_mb_mem[178][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20281_ (.CLK(clknet_leaf_230_clk),
    .D(_01579_),
    .Q(\cur_mb_mem[178][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20282_ (.CLK(clknet_leaf_230_clk),
    .D(_01580_),
    .Q(\cur_mb_mem[178][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20283_ (.CLK(clknet_leaf_50_clk),
    .D(_01581_),
    .Q(\cur_mb_mem[178][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20284_ (.CLK(clknet_leaf_51_clk),
    .D(_01582_),
    .Q(\cur_mb_mem[178][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20285_ (.CLK(clknet_leaf_30_clk),
    .D(_01583_),
    .Q(\cur_mb_mem[179][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20286_ (.CLK(clknet_leaf_42_clk),
    .D(_01584_),
    .Q(\cur_mb_mem[179][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20287_ (.CLK(clknet_leaf_72_clk),
    .D(_01585_),
    .Q(\cur_mb_mem[179][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20288_ (.CLK(clknet_leaf_72_clk),
    .D(_01586_),
    .Q(\cur_mb_mem[179][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20289_ (.CLK(clknet_leaf_356_clk),
    .D(_01587_),
    .Q(\cur_mb_mem[179][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20290_ (.CLK(clknet_leaf_306_clk),
    .D(_01588_),
    .Q(\cur_mb_mem[179][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20291_ (.CLK(clknet_leaf_239_clk),
    .D(_01589_),
    .Q(\cur_mb_mem[179][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20292_ (.CLK(clknet_leaf_46_clk),
    .D(_01590_),
    .Q(\cur_mb_mem[179][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20293_ (.CLK(clknet_leaf_235_clk),
    .D(_01591_),
    .Q(\cur_mb_mem[180][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20294_ (.CLK(clknet_leaf_138_clk),
    .D(_01592_),
    .Q(\cur_mb_mem[180][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20295_ (.CLK(clknet_leaf_235_clk),
    .D(_01593_),
    .Q(\cur_mb_mem[180][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20296_ (.CLK(clknet_leaf_235_clk),
    .D(_01594_),
    .Q(\cur_mb_mem[180][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20297_ (.CLK(clknet_leaf_60_clk),
    .D(_01595_),
    .Q(\cur_mb_mem[180][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20298_ (.CLK(clknet_leaf_57_clk),
    .D(_01596_),
    .Q(\cur_mb_mem[180][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20299_ (.CLK(clknet_leaf_162_clk),
    .D(_01597_),
    .Q(\cur_mb_mem[180][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20300_ (.CLK(clknet_leaf_144_clk),
    .D(_01598_),
    .Q(\cur_mb_mem[180][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20301_ (.CLK(clknet_leaf_349_clk),
    .D(_01599_),
    .Q(\cur_mb_mem[181][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20302_ (.CLK(clknet_leaf_52_clk),
    .D(_01600_),
    .Q(\cur_mb_mem[181][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20303_ (.CLK(clknet_leaf_353_clk),
    .D(_01601_),
    .Q(\cur_mb_mem[181][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20304_ (.CLK(clknet_leaf_352_clk),
    .D(_01602_),
    .Q(\cur_mb_mem[181][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20305_ (.CLK(clknet_leaf_60_clk),
    .D(_01603_),
    .Q(\cur_mb_mem[181][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20306_ (.CLK(clknet_leaf_56_clk),
    .D(_01604_),
    .Q(\cur_mb_mem[181][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20307_ (.CLK(clknet_leaf_355_clk),
    .D(_01605_),
    .Q(\cur_mb_mem[181][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20308_ (.CLK(clknet_leaf_306_clk),
    .D(_01606_),
    .Q(\cur_mb_mem[181][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20309_ (.CLK(clknet_leaf_253_clk),
    .D(_01607_),
    .Q(\cur_mb_mem[182][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20310_ (.CLK(clknet_leaf_238_clk),
    .D(_01608_),
    .Q(\cur_mb_mem[182][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20311_ (.CLK(clknet_leaf_234_clk),
    .D(_01609_),
    .Q(\cur_mb_mem[182][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20312_ (.CLK(clknet_leaf_249_clk),
    .D(_01610_),
    .Q(\cur_mb_mem[182][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20313_ (.CLK(clknet_leaf_232_clk),
    .D(_01611_),
    .Q(\cur_mb_mem[182][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20314_ (.CLK(clknet_leaf_231_clk),
    .D(_01612_),
    .Q(\cur_mb_mem[182][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20315_ (.CLK(clknet_leaf_326_clk),
    .D(_01613_),
    .Q(\cur_mb_mem[182][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20316_ (.CLK(clknet_leaf_325_clk),
    .D(_01614_),
    .Q(\cur_mb_mem[182][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20317_ (.CLK(clknet_leaf_253_clk),
    .D(_01615_),
    .Q(\cur_mb_mem[183][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20318_ (.CLK(clknet_leaf_164_clk),
    .D(_01616_),
    .Q(\cur_mb_mem[183][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20319_ (.CLK(clknet_leaf_234_clk),
    .D(_01617_),
    .Q(\cur_mb_mem[183][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20320_ (.CLK(clknet_leaf_248_clk),
    .D(_01618_),
    .Q(\cur_mb_mem[183][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20321_ (.CLK(clknet_leaf_230_clk),
    .D(_01619_),
    .Q(\cur_mb_mem[183][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20322_ (.CLK(clknet_leaf_230_clk),
    .D(_01620_),
    .Q(\cur_mb_mem[183][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20323_ (.CLK(clknet_leaf_307_clk),
    .D(_01621_),
    .Q(\cur_mb_mem[183][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20324_ (.CLK(clknet_leaf_304_clk),
    .D(_01622_),
    .Q(\cur_mb_mem[183][7] ));
 sky130_fd_sc_hd__dfxtp_2 _20325_ (.CLK(clknet_leaf_341_clk),
    .D(_01623_),
    .Q(\cur_mb_mem[184][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20326_ (.CLK(clknet_leaf_55_clk),
    .D(_01624_),
    .Q(\cur_mb_mem[184][1] ));
 sky130_fd_sc_hd__dfxtp_2 _20327_ (.CLK(clknet_leaf_340_clk),
    .D(_01625_),
    .Q(\cur_mb_mem[184][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20328_ (.CLK(clknet_leaf_341_clk),
    .D(_01626_),
    .Q(\cur_mb_mem[184][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20329_ (.CLK(clknet_leaf_344_clk),
    .D(_01627_),
    .Q(\cur_mb_mem[184][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20330_ (.CLK(clknet_leaf_343_clk),
    .D(_01628_),
    .Q(\cur_mb_mem[184][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20331_ (.CLK(clknet_leaf_51_clk),
    .D(_01629_),
    .Q(\cur_mb_mem[184][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20332_ (.CLK(clknet_leaf_341_clk),
    .D(_01630_),
    .Q(\cur_mb_mem[184][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20333_ (.CLK(clknet_leaf_314_clk),
    .D(_01631_),
    .Q(\cur_mb_mem[185][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20334_ (.CLK(clknet_leaf_307_clk),
    .D(_01632_),
    .Q(\cur_mb_mem[185][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20335_ (.CLK(clknet_leaf_312_clk),
    .D(_01633_),
    .Q(\cur_mb_mem[185][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20336_ (.CLK(clknet_leaf_314_clk),
    .D(_01634_),
    .Q(\cur_mb_mem[185][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20337_ (.CLK(clknet_leaf_344_clk),
    .D(_01635_),
    .Q(\cur_mb_mem[185][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20338_ (.CLK(clknet_leaf_344_clk),
    .D(_01636_),
    .Q(\cur_mb_mem[185][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20339_ (.CLK(clknet_leaf_354_clk),
    .D(_01637_),
    .Q(\cur_mb_mem[185][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20340_ (.CLK(clknet_leaf_354_clk),
    .D(_01638_),
    .Q(\cur_mb_mem[185][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20341_ (.CLK(clknet_leaf_244_clk),
    .D(_01639_),
    .Q(\cur_mb_mem[186][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20342_ (.CLK(clknet_leaf_355_clk),
    .D(_01640_),
    .Q(\cur_mb_mem[186][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20343_ (.CLK(clknet_leaf_43_clk),
    .D(_01641_),
    .Q(\cur_mb_mem[186][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20344_ (.CLK(clknet_leaf_244_clk),
    .D(_01642_),
    .Q(\cur_mb_mem[186][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20345_ (.CLK(clknet_leaf_344_clk),
    .D(_01643_),
    .Q(\cur_mb_mem[186][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20346_ (.CLK(clknet_leaf_343_clk),
    .D(_01644_),
    .Q(\cur_mb_mem[186][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20347_ (.CLK(clknet_leaf_354_clk),
    .D(_01645_),
    .Q(\cur_mb_mem[186][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20348_ (.CLK(clknet_leaf_354_clk),
    .D(_01646_),
    .Q(\cur_mb_mem[186][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20349_ (.CLK(clknet_leaf_308_clk),
    .D(_01647_),
    .Q(\cur_mb_mem[187][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20350_ (.CLK(clknet_leaf_348_clk),
    .D(_01648_),
    .Q(\cur_mb_mem[187][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20351_ (.CLK(clknet_leaf_308_clk),
    .D(_01649_),
    .Q(\cur_mb_mem[187][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20352_ (.CLK(clknet_leaf_306_clk),
    .D(_01650_),
    .Q(\cur_mb_mem[187][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20353_ (.CLK(clknet_leaf_355_clk),
    .D(_01651_),
    .Q(\cur_mb_mem[187][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20354_ (.CLK(clknet_leaf_348_clk),
    .D(_01652_),
    .Q(\cur_mb_mem[187][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20355_ (.CLK(clknet_leaf_307_clk),
    .D(_01653_),
    .Q(\cur_mb_mem[187][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20356_ (.CLK(clknet_leaf_349_clk),
    .D(_01654_),
    .Q(\cur_mb_mem[187][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20357_ (.CLK(clknet_leaf_54_clk),
    .D(_01655_),
    .Q(\cur_mb_mem[188][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20358_ (.CLK(clknet_leaf_54_clk),
    .D(_01656_),
    .Q(\cur_mb_mem[188][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20359_ (.CLK(clknet_leaf_60_clk),
    .D(_01657_),
    .Q(\cur_mb_mem[188][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20360_ (.CLK(clknet_leaf_148_clk),
    .D(_01658_),
    .Q(\cur_mb_mem[188][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20361_ (.CLK(clknet_leaf_356_clk),
    .D(_01659_),
    .Q(\cur_mb_mem[188][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20362_ (.CLK(clknet_leaf_306_clk),
    .D(_01660_),
    .Q(\cur_mb_mem[188][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20363_ (.CLK(clknet_leaf_336_clk),
    .D(_01661_),
    .Q(\cur_mb_mem[188][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20364_ (.CLK(clknet_leaf_324_clk),
    .D(_01662_),
    .Q(\cur_mb_mem[188][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20365_ (.CLK(clknet_leaf_297_clk),
    .D(_01663_),
    .Q(\cur_mb_mem[189][0] ));
 sky130_fd_sc_hd__dfxtp_2 _20366_ (.CLK(clknet_leaf_297_clk),
    .D(_01664_),
    .Q(\cur_mb_mem[189][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20367_ (.CLK(clknet_leaf_299_clk),
    .D(_01665_),
    .Q(\cur_mb_mem[189][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20368_ (.CLK(clknet_leaf_299_clk),
    .D(_01666_),
    .Q(\cur_mb_mem[189][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20369_ (.CLK(clknet_leaf_363_clk),
    .D(_01667_),
    .Q(\cur_mb_mem[189][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20370_ (.CLK(clknet_leaf_299_clk),
    .D(_01668_),
    .Q(\cur_mb_mem[189][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20371_ (.CLK(clknet_leaf_299_clk),
    .D(_01669_),
    .Q(\cur_mb_mem[189][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20372_ (.CLK(clknet_leaf_363_clk),
    .D(_01670_),
    .Q(\cur_mb_mem[189][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20373_ (.CLK(clknet_leaf_388_clk),
    .D(_01671_),
    .Q(\cur_mb_mem[190][0] ));
 sky130_fd_sc_hd__dfxtp_2 _20374_ (.CLK(clknet_leaf_365_clk),
    .D(_01672_),
    .Q(\cur_mb_mem[190][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20375_ (.CLK(clknet_leaf_387_clk),
    .D(_01673_),
    .Q(\cur_mb_mem[190][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20376_ (.CLK(clknet_leaf_389_clk),
    .D(_01674_),
    .Q(\cur_mb_mem[190][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20377_ (.CLK(clknet_leaf_299_clk),
    .D(_01675_),
    .Q(\cur_mb_mem[190][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20378_ (.CLK(clknet_leaf_299_clk),
    .D(_01676_),
    .Q(\cur_mb_mem[190][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20379_ (.CLK(clknet_leaf_370_clk),
    .D(_01677_),
    .Q(\cur_mb_mem[190][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20380_ (.CLK(clknet_leaf_366_clk),
    .D(_01678_),
    .Q(\cur_mb_mem[190][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20381_ (.CLK(clknet_leaf_290_clk),
    .D(_01679_),
    .Q(\cur_mb_mem[191][0] ));
 sky130_fd_sc_hd__dfxtp_2 _20382_ (.CLK(clknet_leaf_297_clk),
    .D(_01680_),
    .Q(\cur_mb_mem[191][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20383_ (.CLK(clknet_leaf_291_clk),
    .D(_01681_),
    .Q(\cur_mb_mem[191][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20384_ (.CLK(clknet_leaf_290_clk),
    .D(_01682_),
    .Q(\cur_mb_mem[191][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20385_ (.CLK(clknet_leaf_297_clk),
    .D(_01683_),
    .Q(\cur_mb_mem[191][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20386_ (.CLK(clknet_leaf_293_clk),
    .D(_01684_),
    .Q(\cur_mb_mem[191][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20387_ (.CLK(clknet_leaf_297_clk),
    .D(_01685_),
    .Q(\cur_mb_mem[191][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20388_ (.CLK(clknet_leaf_298_clk),
    .D(_01686_),
    .Q(\cur_mb_mem[191][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20389_ (.CLK(clknet_leaf_374_clk),
    .D(_01687_),
    .Q(\cur_mb_mem[192][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20390_ (.CLK(clknet_leaf_347_clk),
    .D(_01688_),
    .Q(\cur_mb_mem[192][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20391_ (.CLK(clknet_leaf_53_clk),
    .D(_01689_),
    .Q(\cur_mb_mem[192][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20392_ (.CLK(clknet_leaf_377_clk),
    .D(_01690_),
    .Q(\cur_mb_mem[192][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20393_ (.CLK(clknet_leaf_360_clk),
    .D(_01691_),
    .Q(\cur_mb_mem[192][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20394_ (.CLK(clknet_leaf_360_clk),
    .D(_01692_),
    .Q(\cur_mb_mem[192][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20395_ (.CLK(clknet_leaf_49_clk),
    .D(_01693_),
    .Q(\cur_mb_mem[192][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20396_ (.CLK(clknet_leaf_47_clk),
    .D(_01694_),
    .Q(\cur_mb_mem[192][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20397_ (.CLK(clknet_leaf_8_clk),
    .D(_01695_),
    .Q(\cur_mb_mem[193][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20398_ (.CLK(clknet_leaf_57_clk),
    .D(_01696_),
    .Q(\cur_mb_mem[193][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20399_ (.CLK(clknet_leaf_35_clk),
    .D(_01697_),
    .Q(\cur_mb_mem[193][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20400_ (.CLK(clknet_leaf_10_clk),
    .D(_01698_),
    .Q(\cur_mb_mem[193][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20401_ (.CLK(clknet_leaf_374_clk),
    .D(_01699_),
    .Q(\cur_mb_mem[193][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20402_ (.CLK(clknet_leaf_374_clk),
    .D(_01700_),
    .Q(\cur_mb_mem[193][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20403_ (.CLK(clknet_leaf_346_clk),
    .D(_01701_),
    .Q(\cur_mb_mem[193][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20404_ (.CLK(clknet_leaf_46_clk),
    .D(_01702_),
    .Q(\cur_mb_mem[193][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20405_ (.CLK(clknet_leaf_70_clk),
    .D(_01703_),
    .Q(\cur_mb_mem[194][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20406_ (.CLK(clknet_leaf_238_clk),
    .D(_01704_),
    .Q(\cur_mb_mem[194][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20407_ (.CLK(clknet_leaf_55_clk),
    .D(_01705_),
    .Q(\cur_mb_mem[194][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20408_ (.CLK(clknet_leaf_37_clk),
    .D(_01706_),
    .Q(\cur_mb_mem[194][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20409_ (.CLK(clknet_leaf_375_clk),
    .D(_01707_),
    .Q(\cur_mb_mem[194][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20410_ (.CLK(clknet_leaf_375_clk),
    .D(_01708_),
    .Q(\cur_mb_mem[194][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20411_ (.CLK(clknet_leaf_154_clk),
    .D(_01709_),
    .Q(\cur_mb_mem[194][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20412_ (.CLK(clknet_leaf_238_clk),
    .D(_01710_),
    .Q(\cur_mb_mem[194][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20413_ (.CLK(clknet_leaf_293_clk),
    .D(_01711_),
    .Q(\cur_mb_mem[195][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20414_ (.CLK(clknet_leaf_371_clk),
    .D(_01712_),
    .Q(\cur_mb_mem[195][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20415_ (.CLK(clknet_leaf_293_clk),
    .D(_01713_),
    .Q(\cur_mb_mem[195][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20416_ (.CLK(clknet_leaf_293_clk),
    .D(_01714_),
    .Q(\cur_mb_mem[195][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20417_ (.CLK(clknet_leaf_371_clk),
    .D(_01715_),
    .Q(\cur_mb_mem[195][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20418_ (.CLK(clknet_leaf_370_clk),
    .D(_01716_),
    .Q(\cur_mb_mem[195][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20419_ (.CLK(clknet_leaf_364_clk),
    .D(_01717_),
    .Q(\cur_mb_mem[195][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20420_ (.CLK(clknet_leaf_366_clk),
    .D(_01718_),
    .Q(\cur_mb_mem[195][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20421_ (.CLK(clknet_leaf_383_clk),
    .D(_01719_),
    .Q(\cur_mb_mem[196][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20422_ (.CLK(clknet_leaf_323_clk),
    .D(_01720_),
    .Q(\cur_mb_mem[196][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20423_ (.CLK(clknet_leaf_35_clk),
    .D(_01721_),
    .Q(\cur_mb_mem[196][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20424_ (.CLK(clknet_leaf_383_clk),
    .D(_01722_),
    .Q(\cur_mb_mem[196][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20425_ (.CLK(clknet_leaf_376_clk),
    .D(_01723_),
    .Q(\cur_mb_mem[196][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20426_ (.CLK(clknet_leaf_376_clk),
    .D(_01724_),
    .Q(\cur_mb_mem[196][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20427_ (.CLK(clknet_leaf_40_clk),
    .D(_01725_),
    .Q(\cur_mb_mem[196][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20428_ (.CLK(clknet_leaf_325_clk),
    .D(_01726_),
    .Q(\cur_mb_mem[196][7] ));
 sky130_fd_sc_hd__dfxtp_2 _20429_ (.CLK(clknet_leaf_364_clk),
    .D(_01727_),
    .Q(\cur_mb_mem[197][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20430_ (.CLK(clknet_leaf_371_clk),
    .D(_01728_),
    .Q(\cur_mb_mem[197][1] ));
 sky130_fd_sc_hd__dfxtp_2 _20431_ (.CLK(clknet_leaf_299_clk),
    .D(_01729_),
    .Q(\cur_mb_mem[197][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20432_ (.CLK(clknet_leaf_369_clk),
    .D(_01730_),
    .Q(\cur_mb_mem[197][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20433_ (.CLK(clknet_leaf_387_clk),
    .D(_01731_),
    .Q(\cur_mb_mem[197][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20434_ (.CLK(clknet_leaf_387_clk),
    .D(_01732_),
    .Q(\cur_mb_mem[197][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20435_ (.CLK(clknet_leaf_298_clk),
    .D(_01733_),
    .Q(\cur_mb_mem[197][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20436_ (.CLK(clknet_leaf_363_clk),
    .D(_01734_),
    .Q(\cur_mb_mem[197][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20437_ (.CLK(clknet_leaf_388_clk),
    .D(_01735_),
    .Q(\cur_mb_mem[198][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20438_ (.CLK(clknet_leaf_372_clk),
    .D(_01736_),
    .Q(\cur_mb_mem[198][1] ));
 sky130_fd_sc_hd__dfxtp_2 _20439_ (.CLK(clknet_leaf_387_clk),
    .D(_01737_),
    .Q(\cur_mb_mem[198][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20440_ (.CLK(clknet_leaf_388_clk),
    .D(_01738_),
    .Q(\cur_mb_mem[198][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20441_ (.CLK(clknet_leaf_388_clk),
    .D(_01739_),
    .Q(\cur_mb_mem[198][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20442_ (.CLK(clknet_leaf_388_clk),
    .D(_01740_),
    .Q(\cur_mb_mem[198][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20443_ (.CLK(clknet_leaf_363_clk),
    .D(_01741_),
    .Q(\cur_mb_mem[198][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20444_ (.CLK(clknet_leaf_366_clk),
    .D(_01742_),
    .Q(\cur_mb_mem[198][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20445_ (.CLK(clknet_leaf_291_clk),
    .D(_01743_),
    .Q(\cur_mb_mem[199][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20446_ (.CLK(clknet_leaf_363_clk),
    .D(_01744_),
    .Q(\cur_mb_mem[199][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20447_ (.CLK(clknet_leaf_291_clk),
    .D(_01745_),
    .Q(\cur_mb_mem[199][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20448_ (.CLK(clknet_leaf_292_clk),
    .D(_01746_),
    .Q(\cur_mb_mem[199][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20449_ (.CLK(clknet_leaf_369_clk),
    .D(_01747_),
    .Q(\cur_mb_mem[199][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20450_ (.CLK(clknet_leaf_369_clk),
    .D(_01748_),
    .Q(\cur_mb_mem[199][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20451_ (.CLK(clknet_leaf_297_clk),
    .D(_01749_),
    .Q(\cur_mb_mem[199][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20452_ (.CLK(clknet_leaf_298_clk),
    .D(_01750_),
    .Q(\cur_mb_mem[199][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20453_ (.CLK(clknet_leaf_350_clk),
    .D(_01751_),
    .Q(\cur_mb_mem[200][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20454_ (.CLK(clknet_leaf_45_clk),
    .D(_01752_),
    .Q(\cur_mb_mem[200][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20455_ (.CLK(clknet_leaf_349_clk),
    .D(_01753_),
    .Q(\cur_mb_mem[200][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20456_ (.CLK(clknet_leaf_351_clk),
    .D(_01754_),
    .Q(\cur_mb_mem[200][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20457_ (.CLK(clknet_leaf_376_clk),
    .D(_01755_),
    .Q(\cur_mb_mem[200][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20458_ (.CLK(clknet_leaf_351_clk),
    .D(_01756_),
    .Q(\cur_mb_mem[200][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20459_ (.CLK(clknet_leaf_45_clk),
    .D(_01757_),
    .Q(\cur_mb_mem[200][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20460_ (.CLK(clknet_leaf_48_clk),
    .D(_01758_),
    .Q(\cur_mb_mem[200][7] ));
 sky130_fd_sc_hd__dfxtp_2 _20461_ (.CLK(clknet_leaf_292_clk),
    .D(_01759_),
    .Q(\cur_mb_mem[201][0] ));
 sky130_fd_sc_hd__dfxtp_2 _20462_ (.CLK(clknet_leaf_371_clk),
    .D(_01760_),
    .Q(\cur_mb_mem[201][1] ));
 sky130_fd_sc_hd__dfxtp_2 _20463_ (.CLK(clknet_leaf_292_clk),
    .D(_01761_),
    .Q(\cur_mb_mem[201][2] ));
 sky130_fd_sc_hd__dfxtp_2 _20464_ (.CLK(clknet_leaf_292_clk),
    .D(_01762_),
    .Q(\cur_mb_mem[201][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20465_ (.CLK(clknet_leaf_371_clk),
    .D(_01763_),
    .Q(\cur_mb_mem[201][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20466_ (.CLK(clknet_leaf_370_clk),
    .D(_01764_),
    .Q(\cur_mb_mem[201][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20467_ (.CLK(clknet_leaf_297_clk),
    .D(_01765_),
    .Q(\cur_mb_mem[201][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20468_ (.CLK(clknet_leaf_365_clk),
    .D(_01766_),
    .Q(\cur_mb_mem[201][7] ));
 sky130_fd_sc_hd__dfxtp_2 _20469_ (.CLK(clknet_leaf_372_clk),
    .D(_01767_),
    .Q(\cur_mb_mem[202][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20470_ (.CLK(clknet_leaf_369_clk),
    .D(_01768_),
    .Q(\cur_mb_mem[202][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20471_ (.CLK(clknet_leaf_387_clk),
    .D(_01769_),
    .Q(\cur_mb_mem[202][2] ));
 sky130_fd_sc_hd__dfxtp_2 _20472_ (.CLK(clknet_leaf_372_clk),
    .D(_01770_),
    .Q(\cur_mb_mem[202][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20473_ (.CLK(clknet_leaf_370_clk),
    .D(_01771_),
    .Q(\cur_mb_mem[202][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20474_ (.CLK(clknet_leaf_372_clk),
    .D(_01772_),
    .Q(\cur_mb_mem[202][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20475_ (.CLK(clknet_leaf_365_clk),
    .D(_01773_),
    .Q(\cur_mb_mem[202][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20476_ (.CLK(clknet_leaf_365_clk),
    .D(_01774_),
    .Q(\cur_mb_mem[202][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20477_ (.CLK(clknet_leaf_387_clk),
    .D(_01775_),
    .Q(\cur_mb_mem[203][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20478_ (.CLK(clknet_leaf_372_clk),
    .D(_01776_),
    .Q(\cur_mb_mem[203][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20479_ (.CLK(clknet_leaf_372_clk),
    .D(_01777_),
    .Q(\cur_mb_mem[203][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20480_ (.CLK(clknet_leaf_387_clk),
    .D(_01778_),
    .Q(\cur_mb_mem[203][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20481_ (.CLK(clknet_leaf_366_clk),
    .D(_01779_),
    .Q(\cur_mb_mem[203][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20482_ (.CLK(clknet_leaf_369_clk),
    .D(_01780_),
    .Q(\cur_mb_mem[203][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20483_ (.CLK(clknet_leaf_365_clk),
    .D(_01781_),
    .Q(\cur_mb_mem[203][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20484_ (.CLK(clknet_leaf_365_clk),
    .D(_01782_),
    .Q(\cur_mb_mem[203][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20485_ (.CLK(clknet_leaf_292_clk),
    .D(_01783_),
    .Q(\cur_mb_mem[204][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20486_ (.CLK(clknet_leaf_299_clk),
    .D(_01784_),
    .Q(\cur_mb_mem[204][1] ));
 sky130_fd_sc_hd__dfxtp_2 _20487_ (.CLK(clknet_leaf_295_clk),
    .D(_01785_),
    .Q(\cur_mb_mem[204][2] ));
 sky130_fd_sc_hd__dfxtp_2 _20488_ (.CLK(clknet_leaf_294_clk),
    .D(_01786_),
    .Q(\cur_mb_mem[204][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20489_ (.CLK(clknet_leaf_369_clk),
    .D(_01787_),
    .Q(\cur_mb_mem[204][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20490_ (.CLK(clknet_leaf_369_clk),
    .D(_01788_),
    .Q(\cur_mb_mem[204][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20491_ (.CLK(clknet_leaf_363_clk),
    .D(_01789_),
    .Q(\cur_mb_mem[204][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20492_ (.CLK(clknet_leaf_367_clk),
    .D(_01790_),
    .Q(\cur_mb_mem[204][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20493_ (.CLK(clknet_leaf_372_clk),
    .D(_01791_),
    .Q(\cur_mb_mem[205][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20494_ (.CLK(clknet_leaf_373_clk),
    .D(_01792_),
    .Q(\cur_mb_mem[205][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20495_ (.CLK(clknet_leaf_368_clk),
    .D(_01793_),
    .Q(\cur_mb_mem[205][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20496_ (.CLK(clknet_leaf_373_clk),
    .D(_01794_),
    .Q(\cur_mb_mem[205][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20497_ (.CLK(clknet_leaf_385_clk),
    .D(_01795_),
    .Q(\cur_mb_mem[205][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20498_ (.CLK(clknet_leaf_385_clk),
    .D(_01796_),
    .Q(\cur_mb_mem[205][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20499_ (.CLK(clknet_leaf_368_clk),
    .D(_01797_),
    .Q(\cur_mb_mem[205][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20500_ (.CLK(clknet_leaf_367_clk),
    .D(_01798_),
    .Q(\cur_mb_mem[205][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20501_ (.CLK(clknet_leaf_386_clk),
    .D(_01799_),
    .Q(\cur_mb_mem[206][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20502_ (.CLK(clknet_leaf_372_clk),
    .D(_01800_),
    .Q(\cur_mb_mem[206][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20503_ (.CLK(clknet_leaf_386_clk),
    .D(_01801_),
    .Q(\cur_mb_mem[206][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20504_ (.CLK(clknet_leaf_386_clk),
    .D(_01802_),
    .Q(\cur_mb_mem[206][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20505_ (.CLK(clknet_leaf_361_clk),
    .D(_01803_),
    .Q(\cur_mb_mem[206][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20506_ (.CLK(clknet_leaf_364_clk),
    .D(_01804_),
    .Q(\cur_mb_mem[206][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20507_ (.CLK(clknet_leaf_364_clk),
    .D(_01805_),
    .Q(\cur_mb_mem[206][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20508_ (.CLK(clknet_leaf_363_clk),
    .D(_01806_),
    .Q(\cur_mb_mem[206][7] ));
 sky130_fd_sc_hd__dfxtp_2 _20509_ (.CLK(clknet_leaf_292_clk),
    .D(_01807_),
    .Q(\cur_mb_mem[207][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20510_ (.CLK(clknet_leaf_297_clk),
    .D(_01808_),
    .Q(\cur_mb_mem[207][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20511_ (.CLK(clknet_leaf_294_clk),
    .D(_01809_),
    .Q(\cur_mb_mem[207][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20512_ (.CLK(clknet_leaf_294_clk),
    .D(_01810_),
    .Q(\cur_mb_mem[207][3] ));
 sky130_fd_sc_hd__dfxtp_2 _20513_ (.CLK(clknet_leaf_389_clk),
    .D(_01811_),
    .Q(\cur_mb_mem[207][4] ));
 sky130_fd_sc_hd__dfxtp_2 _20514_ (.CLK(clknet_leaf_386_clk),
    .D(_01812_),
    .Q(\cur_mb_mem[207][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20515_ (.CLK(clknet_leaf_299_clk),
    .D(_01813_),
    .Q(\cur_mb_mem[207][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20516_ (.CLK(clknet_leaf_298_clk),
    .D(_01814_),
    .Q(\cur_mb_mem[207][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20517_ (.CLK(clknet_leaf_383_clk),
    .D(_01815_),
    .Q(\cur_mb_mem[208][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20518_ (.CLK(clknet_leaf_379_clk),
    .D(_01816_),
    .Q(\cur_mb_mem[208][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20519_ (.CLK(clknet_leaf_5_clk),
    .D(_01817_),
    .Q(\cur_mb_mem[208][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20520_ (.CLK(clknet_leaf_383_clk),
    .D(_01818_),
    .Q(\cur_mb_mem[208][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20521_ (.CLK(clknet_leaf_384_clk),
    .D(_01819_),
    .Q(\cur_mb_mem[208][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20522_ (.CLK(clknet_leaf_385_clk),
    .D(_01820_),
    .Q(\cur_mb_mem[208][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20523_ (.CLK(clknet_leaf_358_clk),
    .D(_01821_),
    .Q(\cur_mb_mem[208][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20524_ (.CLK(clknet_leaf_359_clk),
    .D(_01822_),
    .Q(\cur_mb_mem[208][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20525_ (.CLK(clknet_leaf_351_clk),
    .D(_01823_),
    .Q(\cur_mb_mem[209][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20526_ (.CLK(clknet_leaf_354_clk),
    .D(_01824_),
    .Q(\cur_mb_mem[209][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20527_ (.CLK(clknet_leaf_353_clk),
    .D(_01825_),
    .Q(\cur_mb_mem[209][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20528_ (.CLK(clknet_leaf_351_clk),
    .D(_01826_),
    .Q(\cur_mb_mem[209][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20529_ (.CLK(clknet_leaf_358_clk),
    .D(_01827_),
    .Q(\cur_mb_mem[209][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20530_ (.CLK(clknet_leaf_358_clk),
    .D(_01828_),
    .Q(\cur_mb_mem[209][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20531_ (.CLK(clknet_leaf_356_clk),
    .D(_01829_),
    .Q(\cur_mb_mem[209][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20532_ (.CLK(clknet_leaf_358_clk),
    .D(_01830_),
    .Q(\cur_mb_mem[209][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20533_ (.CLK(clknet_leaf_34_clk),
    .D(_01831_),
    .Q(\cur_mb_mem[210][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20534_ (.CLK(clknet_leaf_327_clk),
    .D(_01832_),
    .Q(\cur_mb_mem[210][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20535_ (.CLK(clknet_leaf_32_clk),
    .D(_01833_),
    .Q(\cur_mb_mem[210][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20536_ (.CLK(clknet_leaf_33_clk),
    .D(_01834_),
    .Q(\cur_mb_mem[210][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20537_ (.CLK(clknet_leaf_358_clk),
    .D(_01835_),
    .Q(\cur_mb_mem[210][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20538_ (.CLK(clknet_leaf_352_clk),
    .D(_01836_),
    .Q(\cur_mb_mem[210][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20539_ (.CLK(clknet_leaf_241_clk),
    .D(_01837_),
    .Q(\cur_mb_mem[210][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20540_ (.CLK(clknet_leaf_243_clk),
    .D(_01838_),
    .Q(\cur_mb_mem[210][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20541_ (.CLK(clknet_leaf_389_clk),
    .D(_01839_),
    .Q(\cur_mb_mem[211][0] ));
 sky130_fd_sc_hd__dfxtp_2 _20542_ (.CLK(clknet_leaf_368_clk),
    .D(_01840_),
    .Q(\cur_mb_mem[211][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20543_ (.CLK(clknet_leaf_390_clk),
    .D(_01841_),
    .Q(\cur_mb_mem[211][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20544_ (.CLK(clknet_leaf_390_clk),
    .D(_01842_),
    .Q(\cur_mb_mem[211][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20545_ (.CLK(clknet_leaf_373_clk),
    .D(_01843_),
    .Q(\cur_mb_mem[211][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20546_ (.CLK(clknet_leaf_367_clk),
    .D(_01844_),
    .Q(\cur_mb_mem[211][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20547_ (.CLK(clknet_leaf_370_clk),
    .D(_01845_),
    .Q(\cur_mb_mem[211][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20548_ (.CLK(clknet_leaf_300_clk),
    .D(_01846_),
    .Q(\cur_mb_mem[211][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20549_ (.CLK(clknet_leaf_382_clk),
    .D(_01847_),
    .Q(\cur_mb_mem[212][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20550_ (.CLK(clknet_leaf_348_clk),
    .D(_01848_),
    .Q(\cur_mb_mem[212][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20551_ (.CLK(clknet_leaf_6_clk),
    .D(_01849_),
    .Q(\cur_mb_mem[212][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20552_ (.CLK(clknet_leaf_382_clk),
    .D(_01850_),
    .Q(\cur_mb_mem[212][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20553_ (.CLK(clknet_leaf_383_clk),
    .D(_01851_),
    .Q(\cur_mb_mem[212][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20554_ (.CLK(clknet_leaf_383_clk),
    .D(_01852_),
    .Q(\cur_mb_mem[212][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20555_ (.CLK(clknet_leaf_355_clk),
    .D(_01853_),
    .Q(\cur_mb_mem[212][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20556_ (.CLK(clknet_leaf_357_clk),
    .D(_01854_),
    .Q(\cur_mb_mem[212][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20557_ (.CLK(clknet_leaf_389_clk),
    .D(_01855_),
    .Q(\cur_mb_mem[213][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20558_ (.CLK(clknet_leaf_373_clk),
    .D(_01856_),
    .Q(\cur_mb_mem[213][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20559_ (.CLK(clknet_leaf_390_clk),
    .D(_01857_),
    .Q(\cur_mb_mem[213][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20560_ (.CLK(clknet_leaf_390_clk),
    .D(_01858_),
    .Q(\cur_mb_mem[213][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20561_ (.CLK(clknet_leaf_375_clk),
    .D(_01859_),
    .Q(\cur_mb_mem[213][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20562_ (.CLK(clknet_leaf_368_clk),
    .D(_01860_),
    .Q(\cur_mb_mem[213][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20563_ (.CLK(clknet_leaf_362_clk),
    .D(_01861_),
    .Q(\cur_mb_mem[213][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20564_ (.CLK(clknet_leaf_362_clk),
    .D(_01862_),
    .Q(\cur_mb_mem[213][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20565_ (.CLK(clknet_leaf_293_clk),
    .D(_01863_),
    .Q(\cur_mb_mem[214][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20566_ (.CLK(clknet_leaf_362_clk),
    .D(_01864_),
    .Q(\cur_mb_mem[214][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20567_ (.CLK(clknet_leaf_292_clk),
    .D(_01865_),
    .Q(\cur_mb_mem[214][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20568_ (.CLK(clknet_leaf_294_clk),
    .D(_01866_),
    .Q(\cur_mb_mem[214][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20569_ (.CLK(clknet_leaf_368_clk),
    .D(_01867_),
    .Q(\cur_mb_mem[214][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20570_ (.CLK(clknet_leaf_369_clk),
    .D(_01868_),
    .Q(\cur_mb_mem[214][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20571_ (.CLK(clknet_leaf_364_clk),
    .D(_01869_),
    .Q(\cur_mb_mem[214][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20572_ (.CLK(clknet_leaf_298_clk),
    .D(_01870_),
    .Q(\cur_mb_mem[214][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20573_ (.CLK(clknet_leaf_293_clk),
    .D(_01871_),
    .Q(\cur_mb_mem[215][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20574_ (.CLK(clknet_leaf_363_clk),
    .D(_01872_),
    .Q(\cur_mb_mem[215][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20575_ (.CLK(clknet_leaf_293_clk),
    .D(_01873_),
    .Q(\cur_mb_mem[215][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20576_ (.CLK(clknet_leaf_293_clk),
    .D(_01874_),
    .Q(\cur_mb_mem[215][3] ));
 sky130_fd_sc_hd__dfxtp_2 _20577_ (.CLK(clknet_leaf_371_clk),
    .D(_01875_),
    .Q(\cur_mb_mem[215][4] ));
 sky130_fd_sc_hd__dfxtp_4 _20578_ (.CLK(clknet_leaf_371_clk),
    .D(_01876_),
    .Q(\cur_mb_mem[215][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20579_ (.CLK(clknet_leaf_368_clk),
    .D(_01877_),
    .Q(\cur_mb_mem[215][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20580_ (.CLK(clknet_leaf_364_clk),
    .D(_01878_),
    .Q(\cur_mb_mem[215][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20581_ (.CLK(clknet_leaf_265_clk),
    .D(_01879_),
    .Q(\cur_mb_mem[216][0] ));
 sky130_fd_sc_hd__dfxtp_2 _20582_ (.CLK(clknet_leaf_222_clk),
    .D(_01880_),
    .Q(\cur_mb_mem[216][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20583_ (.CLK(clknet_leaf_265_clk),
    .D(_01881_),
    .Q(\cur_mb_mem[216][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20584_ (.CLK(clknet_leaf_265_clk),
    .D(_01882_),
    .Q(\cur_mb_mem[216][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20585_ (.CLK(clknet_leaf_275_clk),
    .D(_01883_),
    .Q(\cur_mb_mem[216][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20586_ (.CLK(clknet_leaf_275_clk),
    .D(_01884_),
    .Q(\cur_mb_mem[216][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20587_ (.CLK(clknet_leaf_221_clk),
    .D(_01885_),
    .Q(\cur_mb_mem[216][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20588_ (.CLK(clknet_leaf_222_clk),
    .D(_01886_),
    .Q(\cur_mb_mem[216][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20589_ (.CLK(clknet_leaf_389_clk),
    .D(_01887_),
    .Q(\cur_mb_mem[217][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20590_ (.CLK(clknet_leaf_370_clk),
    .D(_01888_),
    .Q(\cur_mb_mem[217][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20591_ (.CLK(clknet_leaf_384_clk),
    .D(_01889_),
    .Q(\cur_mb_mem[217][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20592_ (.CLK(clknet_leaf_389_clk),
    .D(_01890_),
    .Q(\cur_mb_mem[217][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20593_ (.CLK(clknet_leaf_373_clk),
    .D(_01891_),
    .Q(\cur_mb_mem[217][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20594_ (.CLK(clknet_leaf_375_clk),
    .D(_01892_),
    .Q(\cur_mb_mem[217][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20595_ (.CLK(clknet_leaf_300_clk),
    .D(_01893_),
    .Q(\cur_mb_mem[217][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20596_ (.CLK(clknet_leaf_300_clk),
    .D(_01894_),
    .Q(\cur_mb_mem[217][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20597_ (.CLK(clknet_leaf_386_clk),
    .D(_01895_),
    .Q(\cur_mb_mem[218][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20598_ (.CLK(clknet_leaf_373_clk),
    .D(_01896_),
    .Q(\cur_mb_mem[218][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20599_ (.CLK(clknet_leaf_386_clk),
    .D(_01897_),
    .Q(\cur_mb_mem[218][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20600_ (.CLK(clknet_leaf_386_clk),
    .D(_01898_),
    .Q(\cur_mb_mem[218][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20601_ (.CLK(clknet_leaf_362_clk),
    .D(_01899_),
    .Q(\cur_mb_mem[218][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20602_ (.CLK(clknet_leaf_360_clk),
    .D(_01900_),
    .Q(\cur_mb_mem[218][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20603_ (.CLK(clknet_leaf_365_clk),
    .D(_01901_),
    .Q(\cur_mb_mem[218][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20604_ (.CLK(clknet_leaf_367_clk),
    .D(_01902_),
    .Q(\cur_mb_mem[218][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20605_ (.CLK(clknet_leaf_286_clk),
    .D(_01903_),
    .Q(\cur_mb_mem[219][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20606_ (.CLK(clknet_leaf_378_clk),
    .D(_01904_),
    .Q(\cur_mb_mem[219][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20607_ (.CLK(clknet_leaf_312_clk),
    .D(_01905_),
    .Q(\cur_mb_mem[219][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20608_ (.CLK(clknet_leaf_312_clk),
    .D(_01906_),
    .Q(\cur_mb_mem[219][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20609_ (.CLK(clknet_leaf_384_clk),
    .D(_01907_),
    .Q(\cur_mb_mem[219][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20610_ (.CLK(clknet_leaf_381_clk),
    .D(_01908_),
    .Q(\cur_mb_mem[219][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20611_ (.CLK(clknet_leaf_356_clk),
    .D(_01909_),
    .Q(\cur_mb_mem[219][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20612_ (.CLK(clknet_leaf_305_clk),
    .D(_01910_),
    .Q(\cur_mb_mem[219][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20613_ (.CLK(clknet_leaf_384_clk),
    .D(_01911_),
    .Q(\cur_mb_mem[220][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20614_ (.CLK(clknet_leaf_378_clk),
    .D(_01912_),
    .Q(\cur_mb_mem[220][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20615_ (.CLK(clknet_leaf_382_clk),
    .D(_01913_),
    .Q(\cur_mb_mem[220][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20616_ (.CLK(clknet_leaf_382_clk),
    .D(_01914_),
    .Q(\cur_mb_mem[220][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20617_ (.CLK(clknet_leaf_384_clk),
    .D(_01915_),
    .Q(\cur_mb_mem[220][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20618_ (.CLK(clknet_leaf_384_clk),
    .D(_01916_),
    .Q(\cur_mb_mem[220][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20619_ (.CLK(clknet_leaf_305_clk),
    .D(_01917_),
    .Q(\cur_mb_mem[220][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20620_ (.CLK(clknet_leaf_361_clk),
    .D(_01918_),
    .Q(\cur_mb_mem[220][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20621_ (.CLK(clknet_leaf_287_clk),
    .D(_01919_),
    .Q(\cur_mb_mem[221][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20622_ (.CLK(clknet_leaf_376_clk),
    .D(_01920_),
    .Q(\cur_mb_mem[221][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20623_ (.CLK(clknet_leaf_287_clk),
    .D(_01921_),
    .Q(\cur_mb_mem[221][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20624_ (.CLK(clknet_leaf_287_clk),
    .D(_01922_),
    .Q(\cur_mb_mem[221][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20625_ (.CLK(clknet_leaf_385_clk),
    .D(_01923_),
    .Q(\cur_mb_mem[221][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20626_ (.CLK(clknet_leaf_374_clk),
    .D(_01924_),
    .Q(\cur_mb_mem[221][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20627_ (.CLK(clknet_leaf_303_clk),
    .D(_01925_),
    .Q(\cur_mb_mem[221][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20628_ (.CLK(clknet_leaf_360_clk),
    .D(_01926_),
    .Q(\cur_mb_mem[221][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20629_ (.CLK(clknet_leaf_390_clk),
    .D(_01927_),
    .Q(\cur_mb_mem[222][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20630_ (.CLK(clknet_leaf_377_clk),
    .D(_01928_),
    .Q(\cur_mb_mem[222][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20631_ (.CLK(clknet_leaf_382_clk),
    .D(_01929_),
    .Q(\cur_mb_mem[222][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20632_ (.CLK(clknet_leaf_383_clk),
    .D(_01930_),
    .Q(\cur_mb_mem[222][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20633_ (.CLK(clknet_leaf_385_clk),
    .D(_01931_),
    .Q(\cur_mb_mem[222][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20634_ (.CLK(clknet_leaf_374_clk),
    .D(_01932_),
    .Q(\cur_mb_mem[222][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20635_ (.CLK(clknet_leaf_351_clk),
    .D(_01933_),
    .Q(\cur_mb_mem[222][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20636_ (.CLK(clknet_leaf_359_clk),
    .D(_01934_),
    .Q(\cur_mb_mem[222][7] ));
 sky130_fd_sc_hd__dfxtp_2 _20637_ (.CLK(clknet_leaf_295_clk),
    .D(_01935_),
    .Q(\cur_mb_mem[223][0] ));
 sky130_fd_sc_hd__dfxtp_2 _20638_ (.CLK(clknet_leaf_306_clk),
    .D(_01936_),
    .Q(\cur_mb_mem[223][1] ));
 sky130_fd_sc_hd__dfxtp_2 _20639_ (.CLK(clknet_leaf_311_clk),
    .D(_01937_),
    .Q(\cur_mb_mem[223][2] ));
 sky130_fd_sc_hd__dfxtp_2 _20640_ (.CLK(clknet_leaf_311_clk),
    .D(_01938_),
    .Q(\cur_mb_mem[223][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20641_ (.CLK(clknet_leaf_367_clk),
    .D(_01939_),
    .Q(\cur_mb_mem[223][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20642_ (.CLK(clknet_leaf_367_clk),
    .D(_01940_),
    .Q(\cur_mb_mem[223][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20643_ (.CLK(clknet_leaf_310_clk),
    .D(_01941_),
    .Q(\cur_mb_mem[223][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20644_ (.CLK(clknet_leaf_358_clk),
    .D(_01942_),
    .Q(\cur_mb_mem[223][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20645_ (.CLK(clknet_leaf_258_clk),
    .D(_01943_),
    .Q(\cur_mb_mem[224][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20646_ (.CLK(clknet_leaf_259_clk),
    .D(_01944_),
    .Q(\cur_mb_mem[224][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20647_ (.CLK(clknet_leaf_270_clk),
    .D(_01945_),
    .Q(\cur_mb_mem[224][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20648_ (.CLK(clknet_leaf_258_clk),
    .D(_01946_),
    .Q(\cur_mb_mem[224][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20649_ (.CLK(clknet_leaf_280_clk),
    .D(_01947_),
    .Q(\cur_mb_mem[224][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20650_ (.CLK(clknet_leaf_280_clk),
    .D(_01948_),
    .Q(\cur_mb_mem[224][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20651_ (.CLK(clknet_leaf_259_clk),
    .D(_01949_),
    .Q(\cur_mb_mem[224][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20652_ (.CLK(clknet_leaf_303_clk),
    .D(_01950_),
    .Q(\cur_mb_mem[224][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20653_ (.CLK(clknet_leaf_264_clk),
    .D(_01951_),
    .Q(\cur_mb_mem[225][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20654_ (.CLK(clknet_leaf_270_clk),
    .D(_01952_),
    .Q(\cur_mb_mem[225][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20655_ (.CLK(clknet_leaf_223_clk),
    .D(_01953_),
    .Q(\cur_mb_mem[225][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20656_ (.CLK(clknet_leaf_263_clk),
    .D(_01954_),
    .Q(\cur_mb_mem[225][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20657_ (.CLK(clknet_leaf_271_clk),
    .D(_01955_),
    .Q(\cur_mb_mem[225][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20658_ (.CLK(clknet_leaf_272_clk),
    .D(_01956_),
    .Q(\cur_mb_mem[225][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20659_ (.CLK(clknet_leaf_223_clk),
    .D(_01957_),
    .Q(\cur_mb_mem[225][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20660_ (.CLK(clknet_leaf_223_clk),
    .D(_01958_),
    .Q(\cur_mb_mem[225][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20661_ (.CLK(clknet_leaf_269_clk),
    .D(_01959_),
    .Q(\cur_mb_mem[226][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20662_ (.CLK(clknet_leaf_268_clk),
    .D(_01960_),
    .Q(\cur_mb_mem[226][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20663_ (.CLK(clknet_leaf_270_clk),
    .D(_01961_),
    .Q(\cur_mb_mem[226][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20664_ (.CLK(clknet_leaf_269_clk),
    .D(_01962_),
    .Q(\cur_mb_mem[226][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20665_ (.CLK(clknet_leaf_276_clk),
    .D(_01963_),
    .Q(\cur_mb_mem[226][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20666_ (.CLK(clknet_leaf_276_clk),
    .D(_01964_),
    .Q(\cur_mb_mem[226][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20667_ (.CLK(clknet_leaf_268_clk),
    .D(_01965_),
    .Q(\cur_mb_mem[226][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20668_ (.CLK(clknet_leaf_258_clk),
    .D(_01966_),
    .Q(\cur_mb_mem[226][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20669_ (.CLK(clknet_leaf_274_clk),
    .D(_01967_),
    .Q(\cur_mb_mem[227][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20670_ (.CLK(clknet_leaf_314_clk),
    .D(_01968_),
    .Q(\cur_mb_mem[227][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20671_ (.CLK(clknet_leaf_274_clk),
    .D(_01969_),
    .Q(\cur_mb_mem[227][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20672_ (.CLK(clknet_leaf_276_clk),
    .D(_01970_),
    .Q(\cur_mb_mem[227][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20673_ (.CLK(clknet_leaf_276_clk),
    .D(_01971_),
    .Q(\cur_mb_mem[227][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20674_ (.CLK(clknet_leaf_280_clk),
    .D(_01972_),
    .Q(\cur_mb_mem[227][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20675_ (.CLK(clknet_leaf_309_clk),
    .D(_01973_),
    .Q(\cur_mb_mem[227][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20676_ (.CLK(clknet_leaf_304_clk),
    .D(_01974_),
    .Q(\cur_mb_mem[227][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20677_ (.CLK(clknet_5_15__leaf_clk),
    .D(_01975_),
    .Q(\cur_mb_mem[228][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20678_ (.CLK(clknet_leaf_269_clk),
    .D(_01976_),
    .Q(\cur_mb_mem[228][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20679_ (.CLK(clknet_leaf_259_clk),
    .D(_01977_),
    .Q(\cur_mb_mem[228][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20680_ (.CLK(clknet_leaf_269_clk),
    .D(_01978_),
    .Q(\cur_mb_mem[228][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20681_ (.CLK(clknet_leaf_271_clk),
    .D(_01979_),
    .Q(\cur_mb_mem[228][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20682_ (.CLK(clknet_leaf_271_clk),
    .D(_01980_),
    .Q(\cur_mb_mem[228][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20683_ (.CLK(clknet_leaf_265_clk),
    .D(_01981_),
    .Q(\cur_mb_mem[228][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20684_ (.CLK(clknet_leaf_309_clk),
    .D(_01982_),
    .Q(\cur_mb_mem[228][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20685_ (.CLK(clknet_leaf_282_clk),
    .D(_01983_),
    .Q(\cur_mb_mem[229][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20686_ (.CLK(clknet_leaf_283_clk),
    .D(_01984_),
    .Q(\cur_mb_mem[229][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20687_ (.CLK(clknet_leaf_283_clk),
    .D(_01985_),
    .Q(\cur_mb_mem[229][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20688_ (.CLK(clknet_leaf_282_clk),
    .D(_01986_),
    .Q(\cur_mb_mem[229][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20689_ (.CLK(clknet_leaf_284_clk),
    .D(_01987_),
    .Q(\cur_mb_mem[229][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20690_ (.CLK(clknet_leaf_284_clk),
    .D(_01988_),
    .Q(\cur_mb_mem[229][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20691_ (.CLK(clknet_leaf_304_clk),
    .D(_01989_),
    .Q(\cur_mb_mem[229][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20692_ (.CLK(clknet_leaf_304_clk),
    .D(_01990_),
    .Q(\cur_mb_mem[229][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20693_ (.CLK(clknet_leaf_284_clk),
    .D(_01991_),
    .Q(\cur_mb_mem[230][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20694_ (.CLK(clknet_leaf_309_clk),
    .D(_01992_),
    .Q(\cur_mb_mem[230][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20695_ (.CLK(clknet_leaf_285_clk),
    .D(_01993_),
    .Q(\cur_mb_mem[230][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20696_ (.CLK(clknet_leaf_282_clk),
    .D(_01994_),
    .Q(\cur_mb_mem[230][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20697_ (.CLK(clknet_leaf_281_clk),
    .D(_01995_),
    .Q(\cur_mb_mem[230][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20698_ (.CLK(clknet_leaf_281_clk),
    .D(_01996_),
    .Q(\cur_mb_mem[230][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20699_ (.CLK(clknet_leaf_312_clk),
    .D(_01997_),
    .Q(\cur_mb_mem[230][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20700_ (.CLK(clknet_leaf_303_clk),
    .D(_01998_),
    .Q(\cur_mb_mem[230][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20701_ (.CLK(clknet_leaf_275_clk),
    .D(_01999_),
    .Q(\cur_mb_mem[231][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20702_ (.CLK(clknet_leaf_283_clk),
    .D(_02000_),
    .Q(\cur_mb_mem[231][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20703_ (.CLK(clknet_leaf_276_clk),
    .D(_02001_),
    .Q(\cur_mb_mem[231][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20704_ (.CLK(clknet_leaf_274_clk),
    .D(_02002_),
    .Q(\cur_mb_mem[231][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20705_ (.CLK(clknet_leaf_276_clk),
    .D(_02003_),
    .Q(\cur_mb_mem[231][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20706_ (.CLK(clknet_leaf_281_clk),
    .D(_02004_),
    .Q(\cur_mb_mem[231][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20707_ (.CLK(clknet_leaf_312_clk),
    .D(_02005_),
    .Q(\cur_mb_mem[231][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20708_ (.CLK(clknet_leaf_310_clk),
    .D(_02006_),
    .Q(\cur_mb_mem[231][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20709_ (.CLK(clknet_leaf_269_clk),
    .D(_02007_),
    .Q(\cur_mb_mem[232][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20710_ (.CLK(clknet_leaf_268_clk),
    .D(_02008_),
    .Q(\cur_mb_mem[232][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20711_ (.CLK(clknet_leaf_270_clk),
    .D(_02009_),
    .Q(\cur_mb_mem[232][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20712_ (.CLK(clknet_leaf_258_clk),
    .D(_02010_),
    .Q(\cur_mb_mem[232][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20713_ (.CLK(clknet_leaf_276_clk),
    .D(_02011_),
    .Q(\cur_mb_mem[232][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20714_ (.CLK(clknet_leaf_276_clk),
    .D(_02012_),
    .Q(\cur_mb_mem[232][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20715_ (.CLK(clknet_leaf_269_clk),
    .D(_02013_),
    .Q(\cur_mb_mem[232][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20716_ (.CLK(clknet_leaf_258_clk),
    .D(_02014_),
    .Q(\cur_mb_mem[232][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20717_ (.CLK(clknet_leaf_284_clk),
    .D(_02015_),
    .Q(\cur_mb_mem[233][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20718_ (.CLK(clknet_leaf_284_clk),
    .D(_02016_),
    .Q(\cur_mb_mem[233][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20719_ (.CLK(clknet_leaf_284_clk),
    .D(_02017_),
    .Q(\cur_mb_mem[233][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20720_ (.CLK(clknet_leaf_285_clk),
    .D(_02018_),
    .Q(\cur_mb_mem[233][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20721_ (.CLK(clknet_leaf_281_clk),
    .D(_02019_),
    .Q(\cur_mb_mem[233][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20722_ (.CLK(clknet_leaf_281_clk),
    .D(_02020_),
    .Q(\cur_mb_mem[233][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20723_ (.CLK(clknet_leaf_310_clk),
    .D(_02021_),
    .Q(\cur_mb_mem[233][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20724_ (.CLK(clknet_leaf_310_clk),
    .D(_02022_),
    .Q(\cur_mb_mem[233][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20725_ (.CLK(clknet_leaf_277_clk),
    .D(_02023_),
    .Q(\cur_mb_mem[234][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20726_ (.CLK(clknet_leaf_295_clk),
    .D(_02024_),
    .Q(\cur_mb_mem[234][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20727_ (.CLK(clknet_leaf_279_clk),
    .D(_02025_),
    .Q(\cur_mb_mem[234][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20728_ (.CLK(clknet_leaf_277_clk),
    .D(_02026_),
    .Q(\cur_mb_mem[234][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20729_ (.CLK(clknet_leaf_279_clk),
    .D(_02027_),
    .Q(\cur_mb_mem[234][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20730_ (.CLK(clknet_leaf_279_clk),
    .D(_02028_),
    .Q(\cur_mb_mem[234][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20731_ (.CLK(clknet_leaf_295_clk),
    .D(_02029_),
    .Q(\cur_mb_mem[234][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20732_ (.CLK(clknet_leaf_302_clk),
    .D(_02030_),
    .Q(\cur_mb_mem[234][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20733_ (.CLK(clknet_leaf_277_clk),
    .D(_02031_),
    .Q(\cur_mb_mem[235][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20734_ (.CLK(clknet_leaf_289_clk),
    .D(_02032_),
    .Q(\cur_mb_mem[235][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20735_ (.CLK(clknet_leaf_277_clk),
    .D(_02033_),
    .Q(\cur_mb_mem[235][2] ));
 sky130_fd_sc_hd__dfxtp_2 _20736_ (.CLK(clknet_leaf_277_clk),
    .D(_02034_),
    .Q(\cur_mb_mem[235][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20737_ (.CLK(clknet_leaf_278_clk),
    .D(_02035_),
    .Q(\cur_mb_mem[235][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20738_ (.CLK(clknet_leaf_278_clk),
    .D(_02036_),
    .Q(\cur_mb_mem[235][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20739_ (.CLK(clknet_leaf_295_clk),
    .D(_02037_),
    .Q(\cur_mb_mem[235][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20740_ (.CLK(clknet_leaf_296_clk),
    .D(_02038_),
    .Q(\cur_mb_mem[235][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20741_ (.CLK(clknet_leaf_285_clk),
    .D(_02039_),
    .Q(\cur_mb_mem[236][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20742_ (.CLK(clknet_leaf_285_clk),
    .D(_02040_),
    .Q(\cur_mb_mem[236][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20743_ (.CLK(clknet_leaf_277_clk),
    .D(_02041_),
    .Q(\cur_mb_mem[236][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20744_ (.CLK(clknet_leaf_288_clk),
    .D(_02042_),
    .Q(\cur_mb_mem[236][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20745_ (.CLK(clknet_leaf_278_clk),
    .D(_02043_),
    .Q(\cur_mb_mem[236][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20746_ (.CLK(clknet_leaf_281_clk),
    .D(_02044_),
    .Q(\cur_mb_mem[236][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20747_ (.CLK(clknet_leaf_295_clk),
    .D(_02045_),
    .Q(\cur_mb_mem[236][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20748_ (.CLK(clknet_leaf_302_clk),
    .D(_02046_),
    .Q(\cur_mb_mem[236][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20749_ (.CLK(clknet_leaf_286_clk),
    .D(_02047_),
    .Q(\cur_mb_mem[237][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20750_ (.CLK(clknet_leaf_289_clk),
    .D(_02048_),
    .Q(\cur_mb_mem[237][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20751_ (.CLK(clknet_leaf_294_clk),
    .D(_02049_),
    .Q(\cur_mb_mem[237][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20752_ (.CLK(clknet_leaf_292_clk),
    .D(_02050_),
    .Q(\cur_mb_mem[237][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20753_ (.CLK(clknet_leaf_288_clk),
    .D(_02051_),
    .Q(\cur_mb_mem[237][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20754_ (.CLK(clknet_leaf_288_clk),
    .D(_02052_),
    .Q(\cur_mb_mem[237][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20755_ (.CLK(clknet_leaf_296_clk),
    .D(_02053_),
    .Q(\cur_mb_mem[237][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20756_ (.CLK(clknet_leaf_296_clk),
    .D(_02054_),
    .Q(\cur_mb_mem[237][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20757_ (.CLK(clknet_leaf_295_clk),
    .D(_02055_),
    .Q(\cur_mb_mem[238][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20758_ (.CLK(clknet_leaf_287_clk),
    .D(_02056_),
    .Q(\cur_mb_mem[238][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20759_ (.CLK(clknet_leaf_361_clk),
    .D(_02057_),
    .Q(\cur_mb_mem[238][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20760_ (.CLK(clknet_leaf_294_clk),
    .D(_02058_),
    .Q(\cur_mb_mem[238][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20761_ (.CLK(clknet_leaf_361_clk),
    .D(_02059_),
    .Q(\cur_mb_mem[238][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20762_ (.CLK(clknet_leaf_361_clk),
    .D(_02060_),
    .Q(\cur_mb_mem[238][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20763_ (.CLK(clknet_leaf_300_clk),
    .D(_02061_),
    .Q(\cur_mb_mem[238][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20764_ (.CLK(clknet_leaf_302_clk),
    .D(_02062_),
    .Q(\cur_mb_mem[238][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20765_ (.CLK(clknet_leaf_289_clk),
    .D(_02063_),
    .Q(\cur_mb_mem[239][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20766_ (.CLK(clknet_leaf_289_clk),
    .D(_02064_),
    .Q(\cur_mb_mem[239][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20767_ (.CLK(clknet_leaf_290_clk),
    .D(_02065_),
    .Q(\cur_mb_mem[239][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20768_ (.CLK(clknet_leaf_289_clk),
    .D(_02066_),
    .Q(\cur_mb_mem[239][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20769_ (.CLK(clknet_leaf_287_clk),
    .D(_02067_),
    .Q(\cur_mb_mem[239][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20770_ (.CLK(clknet_leaf_287_clk),
    .D(_02068_),
    .Q(\cur_mb_mem[239][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20771_ (.CLK(clknet_leaf_296_clk),
    .D(_02069_),
    .Q(\cur_mb_mem[239][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20772_ (.CLK(clknet_leaf_296_clk),
    .D(_02070_),
    .Q(\cur_mb_mem[239][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20773_ (.CLK(clknet_leaf_269_clk),
    .D(_02071_),
    .Q(\cur_mb_mem[240][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20774_ (.CLK(clknet_leaf_268_clk),
    .D(_02072_),
    .Q(\cur_mb_mem[240][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20775_ (.CLK(clknet_leaf_223_clk),
    .D(_02073_),
    .Q(\cur_mb_mem[240][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20776_ (.CLK(clknet_leaf_264_clk),
    .D(_02074_),
    .Q(\cur_mb_mem[240][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20777_ (.CLK(clknet_leaf_275_clk),
    .D(_02075_),
    .Q(\cur_mb_mem[240][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20778_ (.CLK(clknet_leaf_275_clk),
    .D(_02076_),
    .Q(\cur_mb_mem[240][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20779_ (.CLK(clknet_leaf_259_clk),
    .D(_02077_),
    .Q(\cur_mb_mem[240][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20780_ (.CLK(clknet_leaf_223_clk),
    .D(_02078_),
    .Q(\cur_mb_mem[240][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20781_ (.CLK(clknet_leaf_259_clk),
    .D(_02079_),
    .Q(\cur_mb_mem[241][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20782_ (.CLK(clknet_leaf_271_clk),
    .D(_02080_),
    .Q(\cur_mb_mem[241][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20783_ (.CLK(clknet_leaf_222_clk),
    .D(_02081_),
    .Q(\cur_mb_mem[241][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20784_ (.CLK(clknet_leaf_260_clk),
    .D(_02082_),
    .Q(\cur_mb_mem[241][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20785_ (.CLK(clknet_leaf_276_clk),
    .D(_02083_),
    .Q(\cur_mb_mem[241][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20786_ (.CLK(clknet_leaf_276_clk),
    .D(_02084_),
    .Q(\cur_mb_mem[241][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20787_ (.CLK(clknet_leaf_259_clk),
    .D(_02085_),
    .Q(\cur_mb_mem[241][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20788_ (.CLK(clknet_leaf_260_clk),
    .D(_02086_),
    .Q(\cur_mb_mem[241][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20789_ (.CLK(clknet_leaf_265_clk),
    .D(_02087_),
    .Q(\cur_mb_mem[242][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20790_ (.CLK(clknet_leaf_222_clk),
    .D(_02088_),
    .Q(\cur_mb_mem[242][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20791_ (.CLK(clknet_leaf_264_clk),
    .D(_02089_),
    .Q(\cur_mb_mem[242][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20792_ (.CLK(clknet_5_15__leaf_clk),
    .D(_02090_),
    .Q(\cur_mb_mem[242][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20793_ (.CLK(clknet_leaf_271_clk),
    .D(_02091_),
    .Q(\cur_mb_mem[242][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20794_ (.CLK(clknet_leaf_268_clk),
    .D(_02092_),
    .Q(\cur_mb_mem[242][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20795_ (.CLK(clknet_leaf_264_clk),
    .D(_02093_),
    .Q(\cur_mb_mem[242][6] ));
 sky130_fd_sc_hd__dfxtp_2 _20796_ (.CLK(clknet_leaf_264_clk),
    .D(_02094_),
    .Q(\cur_mb_mem[242][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20797_ (.CLK(clknet_leaf_278_clk),
    .D(_02095_),
    .Q(\cur_mb_mem[243][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20798_ (.CLK(clknet_leaf_289_clk),
    .D(_02096_),
    .Q(\cur_mb_mem[243][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20799_ (.CLK(clknet_leaf_289_clk),
    .D(_02097_),
    .Q(\cur_mb_mem[243][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20800_ (.CLK(clknet_leaf_277_clk),
    .D(_02098_),
    .Q(\cur_mb_mem[243][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20801_ (.CLK(clknet_leaf_280_clk),
    .D(_02099_),
    .Q(\cur_mb_mem[243][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20802_ (.CLK(clknet_leaf_280_clk),
    .D(_02100_),
    .Q(\cur_mb_mem[243][5] ));
 sky130_fd_sc_hd__dfxtp_2 _20803_ (.CLK(clknet_leaf_300_clk),
    .D(_02101_),
    .Q(\cur_mb_mem[243][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20804_ (.CLK(clknet_leaf_301_clk),
    .D(_02102_),
    .Q(\cur_mb_mem[243][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20805_ (.CLK(clknet_leaf_263_clk),
    .D(_02103_),
    .Q(\cur_mb_mem[244][0] ));
 sky130_fd_sc_hd__dfxtp_4 _20806_ (.CLK(clknet_leaf_224_clk),
    .D(_02104_),
    .Q(\cur_mb_mem[244][1] ));
 sky130_fd_sc_hd__dfxtp_2 _20807_ (.CLK(clknet_leaf_222_clk),
    .D(_02105_),
    .Q(\cur_mb_mem[244][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20808_ (.CLK(clknet_leaf_263_clk),
    .D(_02106_),
    .Q(\cur_mb_mem[244][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20809_ (.CLK(clknet_leaf_295_clk),
    .D(_02107_),
    .Q(\cur_mb_mem[244][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20810_ (.CLK(clknet_leaf_295_clk),
    .D(_02108_),
    .Q(\cur_mb_mem[244][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20811_ (.CLK(clknet_leaf_257_clk),
    .D(_02109_),
    .Q(\cur_mb_mem[244][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20812_ (.CLK(clknet_leaf_295_clk),
    .D(_02110_),
    .Q(\cur_mb_mem[244][7] ));
 sky130_fd_sc_hd__dfxtp_4 _20813_ (.CLK(clknet_leaf_302_clk),
    .D(_02111_),
    .Q(\cur_mb_mem[245][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20814_ (.CLK(clknet_leaf_301_clk),
    .D(_02112_),
    .Q(\cur_mb_mem[245][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20815_ (.CLK(clknet_leaf_367_clk),
    .D(_02113_),
    .Q(\cur_mb_mem[245][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20816_ (.CLK(clknet_leaf_302_clk),
    .D(_02114_),
    .Q(\cur_mb_mem[245][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20817_ (.CLK(clknet_leaf_367_clk),
    .D(_02115_),
    .Q(\cur_mb_mem[245][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20818_ (.CLK(clknet_leaf_367_clk),
    .D(_02116_),
    .Q(\cur_mb_mem[245][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20819_ (.CLK(clknet_leaf_301_clk),
    .D(_02117_),
    .Q(\cur_mb_mem[245][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20820_ (.CLK(clknet_leaf_301_clk),
    .D(_02118_),
    .Q(\cur_mb_mem[245][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20821_ (.CLK(clknet_leaf_278_clk),
    .D(_02119_),
    .Q(\cur_mb_mem[246][0] ));
 sky130_fd_sc_hd__dfxtp_2 _20822_ (.CLK(clknet_leaf_361_clk),
    .D(_02120_),
    .Q(\cur_mb_mem[246][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20823_ (.CLK(clknet_leaf_289_clk),
    .D(_02121_),
    .Q(\cur_mb_mem[246][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20824_ (.CLK(clknet_leaf_277_clk),
    .D(_02122_),
    .Q(\cur_mb_mem[246][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20825_ (.CLK(clknet_leaf_279_clk),
    .D(_02123_),
    .Q(\cur_mb_mem[246][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20826_ (.CLK(clknet_leaf_279_clk),
    .D(_02124_),
    .Q(\cur_mb_mem[246][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20827_ (.CLK(clknet_leaf_361_clk),
    .D(_02125_),
    .Q(\cur_mb_mem[246][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20828_ (.CLK(clknet_leaf_301_clk),
    .D(_02126_),
    .Q(\cur_mb_mem[246][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20829_ (.CLK(clknet_leaf_288_clk),
    .D(_02127_),
    .Q(\cur_mb_mem[247][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20830_ (.CLK(clknet_leaf_367_clk),
    .D(_02128_),
    .Q(\cur_mb_mem[247][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20831_ (.CLK(clknet_leaf_294_clk),
    .D(_02129_),
    .Q(\cur_mb_mem[247][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20832_ (.CLK(clknet_leaf_288_clk),
    .D(_02130_),
    .Q(\cur_mb_mem[247][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20833_ (.CLK(clknet_leaf_359_clk),
    .D(_02131_),
    .Q(\cur_mb_mem[247][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20834_ (.CLK(clknet_leaf_359_clk),
    .D(_02132_),
    .Q(\cur_mb_mem[247][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20835_ (.CLK(clknet_leaf_296_clk),
    .D(_02133_),
    .Q(\cur_mb_mem[247][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20836_ (.CLK(clknet_leaf_298_clk),
    .D(_02134_),
    .Q(\cur_mb_mem[247][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20837_ (.CLK(clknet_leaf_314_clk),
    .D(_02135_),
    .Q(\cur_mb_mem[248][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20838_ (.CLK(clknet_leaf_224_clk),
    .D(_02136_),
    .Q(\cur_mb_mem[248][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20839_ (.CLK(clknet_leaf_283_clk),
    .D(_02137_),
    .Q(\cur_mb_mem[248][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20840_ (.CLK(clknet_leaf_261_clk),
    .D(_02138_),
    .Q(\cur_mb_mem[248][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20841_ (.CLK(clknet_leaf_274_clk),
    .D(_02139_),
    .Q(\cur_mb_mem[248][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20842_ (.CLK(clknet_leaf_274_clk),
    .D(_02140_),
    .Q(\cur_mb_mem[248][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20843_ (.CLK(clknet_leaf_235_clk),
    .D(_02141_),
    .Q(\cur_mb_mem[248][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20844_ (.CLK(clknet_leaf_319_clk),
    .D(_02142_),
    .Q(\cur_mb_mem[248][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20845_ (.CLK(clknet_leaf_4_clk),
    .D(_02143_),
    .Q(\cur_mb_mem[249][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20846_ (.CLK(clknet_leaf_344_clk),
    .D(_02144_),
    .Q(\cur_mb_mem[249][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20847_ (.CLK(clknet_leaf_5_clk),
    .D(_02145_),
    .Q(\cur_mb_mem[249][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20848_ (.CLK(clknet_leaf_4_clk),
    .D(_02146_),
    .Q(\cur_mb_mem[249][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20849_ (.CLK(clknet_leaf_282_clk),
    .D(_02147_),
    .Q(\cur_mb_mem[249][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20850_ (.CLK(clknet_leaf_282_clk),
    .D(_02148_),
    .Q(\cur_mb_mem[249][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20851_ (.CLK(clknet_leaf_337_clk),
    .D(_02149_),
    .Q(\cur_mb_mem[249][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20852_ (.CLK(clknet_leaf_342_clk),
    .D(_02150_),
    .Q(\cur_mb_mem[249][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20853_ (.CLK(clknet_leaf_4_clk),
    .D(_02151_),
    .Q(\cur_mb_mem[250][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20854_ (.CLK(clknet_leaf_342_clk),
    .D(_02152_),
    .Q(\cur_mb_mem[250][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20855_ (.CLK(clknet_leaf_5_clk),
    .D(_02153_),
    .Q(\cur_mb_mem[250][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20856_ (.CLK(clknet_leaf_4_clk),
    .D(_02154_),
    .Q(\cur_mb_mem[250][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20857_ (.CLK(clknet_leaf_383_clk),
    .D(_02155_),
    .Q(\cur_mb_mem[250][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20858_ (.CLK(clknet_leaf_384_clk),
    .D(_02156_),
    .Q(\cur_mb_mem[250][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20859_ (.CLK(clknet_leaf_358_clk),
    .D(_02157_),
    .Q(\cur_mb_mem[250][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20860_ (.CLK(clknet_leaf_341_clk),
    .D(_02158_),
    .Q(\cur_mb_mem[250][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20861_ (.CLK(clknet_leaf_35_clk),
    .D(_02159_),
    .Q(\cur_mb_mem[251][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20862_ (.CLK(clknet_leaf_40_clk),
    .D(_02160_),
    .Q(\cur_mb_mem[251][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20863_ (.CLK(clknet_leaf_34_clk),
    .D(_02161_),
    .Q(\cur_mb_mem[251][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20864_ (.CLK(clknet_leaf_35_clk),
    .D(_02162_),
    .Q(\cur_mb_mem[251][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20865_ (.CLK(clknet_leaf_272_clk),
    .D(_02163_),
    .Q(\cur_mb_mem[251][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20866_ (.CLK(clknet_leaf_271_clk),
    .D(_02164_),
    .Q(\cur_mb_mem[251][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20867_ (.CLK(clknet_leaf_40_clk),
    .D(_02165_),
    .Q(\cur_mb_mem[251][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20868_ (.CLK(clknet_leaf_342_clk),
    .D(_02166_),
    .Q(\cur_mb_mem[251][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20869_ (.CLK(clknet_leaf_32_clk),
    .D(_02167_),
    .Q(\cur_mb_mem[252][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20870_ (.CLK(clknet_leaf_346_clk),
    .D(_02168_),
    .Q(\cur_mb_mem[252][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20871_ (.CLK(clknet_leaf_31_clk),
    .D(_02169_),
    .Q(\cur_mb_mem[252][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20872_ (.CLK(clknet_leaf_32_clk),
    .D(_02170_),
    .Q(\cur_mb_mem[252][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20873_ (.CLK(clknet_leaf_377_clk),
    .D(_02171_),
    .Q(\cur_mb_mem[252][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20874_ (.CLK(clknet_leaf_378_clk),
    .D(_02172_),
    .Q(\cur_mb_mem[252][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20875_ (.CLK(clknet_leaf_336_clk),
    .D(_02173_),
    .Q(\cur_mb_mem[252][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20876_ (.CLK(clknet_leaf_357_clk),
    .D(_02174_),
    .Q(\cur_mb_mem[252][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20877_ (.CLK(clknet_leaf_380_clk),
    .D(_02175_),
    .Q(\cur_mb_mem[253][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20878_ (.CLK(clknet_leaf_346_clk),
    .D(_02176_),
    .Q(\cur_mb_mem[253][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20879_ (.CLK(clknet_leaf_6_clk),
    .D(_02177_),
    .Q(\cur_mb_mem[253][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20880_ (.CLK(clknet_leaf_381_clk),
    .D(_02178_),
    .Q(\cur_mb_mem[253][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20881_ (.CLK(clknet_leaf_375_clk),
    .D(_02179_),
    .Q(\cur_mb_mem[253][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20882_ (.CLK(clknet_leaf_374_clk),
    .D(_02180_),
    .Q(\cur_mb_mem[253][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20883_ (.CLK(clknet_leaf_340_clk),
    .D(_02181_),
    .Q(\cur_mb_mem[253][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20884_ (.CLK(clknet_leaf_340_clk),
    .D(_02182_),
    .Q(\cur_mb_mem[253][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20885_ (.CLK(clknet_leaf_6_clk),
    .D(_02183_),
    .Q(\cur_mb_mem[254][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20886_ (.CLK(clknet_leaf_354_clk),
    .D(_02184_),
    .Q(\cur_mb_mem[254][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20887_ (.CLK(clknet_leaf_6_clk),
    .D(_02185_),
    .Q(\cur_mb_mem[254][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20888_ (.CLK(clknet_leaf_381_clk),
    .D(_02186_),
    .Q(\cur_mb_mem[254][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20889_ (.CLK(clknet_leaf_275_clk),
    .D(_02187_),
    .Q(\cur_mb_mem[254][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20890_ (.CLK(clknet_leaf_275_clk),
    .D(_02188_),
    .Q(\cur_mb_mem[254][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20891_ (.CLK(clknet_leaf_357_clk),
    .D(_02189_),
    .Q(\cur_mb_mem[254][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20892_ (.CLK(clknet_leaf_358_clk),
    .D(_02190_),
    .Q(\cur_mb_mem[254][7] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9179 ();
 sky130_fd_sc_hd__buf_4 input1 (.A(frame_start_addr[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input2 (.A(frame_start_addr[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(frame_start_addr[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(frame_start_addr[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_6 input5 (.A(frame_start_addr[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(frame_start_addr[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(frame_start_addr[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(frame_start_addr[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(frame_start_addr[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input10 (.A(frame_start_addr[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(frame_start_addr[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_8 input12 (.A(frame_start_addr[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(frame_start_addr[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_8 input14 (.A(frame_start_addr[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(frame_start_addr[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_8 input16 (.A(frame_start_addr[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(frame_start_addr[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(frame_start_addr[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_6 input19 (.A(frame_start_addr[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(frame_start_addr[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(frame_start_addr[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(frame_start_addr[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(frame_start_addr[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_8 input24 (.A(frame_start_addr[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(frame_start_addr[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(frame_start_addr[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(frame_start_addr[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(frame_start_addr[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(frame_start_addr[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(frame_start_addr[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(frame_start_addr[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(frame_start_addr[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(mb_x_pos[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(mb_x_pos[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(mb_x_pos[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_6 input36 (.A(mb_x_pos[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(mb_x_pos[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(mb_x_pos[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_6 input39 (.A(mb_x_pos[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_8 input40 (.A(mb_x_pos[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_8 input41 (.A(mb_x_pos[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_8 input42 (.A(mb_x_pos[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(mb_x_pos[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_4 input44 (.A(mb_x_pos[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_4 input45 (.A(mb_x_pos[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_16 input46 (.A(mb_x_pos[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_6 input47 (.A(mb_x_pos[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(mb_x_pos[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_8 input49 (.A(mb_x_pos[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_8 input50 (.A(mb_x_pos[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input51 (.A(mb_x_pos[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_8 input52 (.A(mb_x_pos[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(mb_x_pos[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_8 input54 (.A(mb_x_pos[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_4 input55 (.A(mb_x_pos[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_6 input56 (.A(mb_x_pos[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_8 input57 (.A(mb_x_pos[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_8 input58 (.A(mb_x_pos[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_8 input59 (.A(mb_x_pos[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_8 input60 (.A(mb_x_pos[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 input61 (.A(mb_x_pos[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_8 input62 (.A(mb_x_pos[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_8 input63 (.A(mb_x_pos[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(mb_x_pos[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(mb_y_pos[0]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_16 input66 (.A(mb_y_pos[10]),
    .X(net66));
 sky130_fd_sc_hd__buf_2 input67 (.A(mb_y_pos[11]),
    .X(net67));
 sky130_fd_sc_hd__buf_8 input68 (.A(mb_y_pos[12]),
    .X(net68));
 sky130_fd_sc_hd__buf_4 input69 (.A(mb_y_pos[13]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_16 input70 (.A(mb_y_pos[14]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_8 input71 (.A(mb_y_pos[15]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 input72 (.A(mb_y_pos[16]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(mb_y_pos[17]),
    .X(net73));
 sky130_fd_sc_hd__buf_4 input74 (.A(mb_y_pos[18]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 input75 (.A(mb_y_pos[19]),
    .X(net75));
 sky130_fd_sc_hd__buf_6 input76 (.A(mb_y_pos[1]),
    .X(net76));
 sky130_fd_sc_hd__buf_4 input77 (.A(mb_y_pos[20]),
    .X(net77));
 sky130_fd_sc_hd__buf_8 input78 (.A(mb_y_pos[21]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 input79 (.A(mb_y_pos[22]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_16 input80 (.A(mb_y_pos[23]),
    .X(net80));
 sky130_fd_sc_hd__buf_2 input81 (.A(mb_y_pos[24]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(mb_y_pos[25]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_8 input83 (.A(mb_y_pos[26]),
    .X(net83));
 sky130_fd_sc_hd__buf_8 input84 (.A(mb_y_pos[27]),
    .X(net84));
 sky130_fd_sc_hd__buf_6 input85 (.A(mb_y_pos[28]),
    .X(net85));
 sky130_fd_sc_hd__buf_8 input86 (.A(mb_y_pos[29]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(mb_y_pos[2]),
    .X(net87));
 sky130_fd_sc_hd__buf_2 input88 (.A(mb_y_pos[30]),
    .X(net88));
 sky130_fd_sc_hd__buf_6 input89 (.A(mb_y_pos[31]),
    .X(net89));
 sky130_fd_sc_hd__buf_6 input90 (.A(mb_y_pos[3]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 input91 (.A(mb_y_pos[4]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_8 input92 (.A(mb_y_pos[5]),
    .X(net92));
 sky130_fd_sc_hd__buf_8 input93 (.A(mb_y_pos[6]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(mb_y_pos[7]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 input95 (.A(mb_y_pos[8]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_8 input96 (.A(mb_y_pos[9]),
    .X(net96));
 sky130_fd_sc_hd__buf_12 input97 (.A(mem_rdata[0]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_16 input98 (.A(mem_rdata[1]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_16 input99 (.A(mem_rdata[2]),
    .X(net99));
 sky130_fd_sc_hd__buf_12 input100 (.A(mem_rdata[3]),
    .X(net100));
 sky130_fd_sc_hd__buf_12 input101 (.A(mem_rdata[4]),
    .X(net101));
 sky130_fd_sc_hd__buf_12 input102 (.A(mem_rdata[5]),
    .X(net102));
 sky130_fd_sc_hd__buf_12 input103 (.A(mem_rdata[6]),
    .X(net103));
 sky130_fd_sc_hd__buf_8 input104 (.A(mem_rdata[7]),
    .X(net104));
 sky130_fd_sc_hd__buf_6 input105 (.A(ref_start_addr[0]),
    .X(net105));
 sky130_fd_sc_hd__buf_2 input106 (.A(ref_start_addr[10]),
    .X(net106));
 sky130_fd_sc_hd__buf_4 input107 (.A(ref_start_addr[11]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 input108 (.A(ref_start_addr[12]),
    .X(net108));
 sky130_fd_sc_hd__buf_8 input109 (.A(ref_start_addr[13]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 input110 (.A(ref_start_addr[14]),
    .X(net110));
 sky130_fd_sc_hd__buf_6 input111 (.A(ref_start_addr[15]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_8 input112 (.A(ref_start_addr[16]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(ref_start_addr[17]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 input114 (.A(ref_start_addr[18]),
    .X(net114));
 sky130_fd_sc_hd__buf_2 input115 (.A(ref_start_addr[19]),
    .X(net115));
 sky130_fd_sc_hd__buf_4 input116 (.A(ref_start_addr[1]),
    .X(net116));
 sky130_fd_sc_hd__buf_6 input117 (.A(ref_start_addr[20]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(ref_start_addr[21]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_8 input119 (.A(ref_start_addr[22]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input120 (.A(ref_start_addr[23]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 input121 (.A(ref_start_addr[24]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 input122 (.A(ref_start_addr[25]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 input123 (.A(ref_start_addr[26]),
    .X(net123));
 sky130_fd_sc_hd__buf_6 input124 (.A(ref_start_addr[27]),
    .X(net124));
 sky130_fd_sc_hd__buf_6 input125 (.A(ref_start_addr[28]),
    .X(net125));
 sky130_fd_sc_hd__buf_4 input126 (.A(ref_start_addr[29]),
    .X(net126));
 sky130_fd_sc_hd__buf_8 input127 (.A(ref_start_addr[2]),
    .X(net127));
 sky130_fd_sc_hd__buf_6 input128 (.A(ref_start_addr[30]),
    .X(net128));
 sky130_fd_sc_hd__buf_6 input129 (.A(ref_start_addr[31]),
    .X(net129));
 sky130_fd_sc_hd__buf_4 input130 (.A(ref_start_addr[3]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(ref_start_addr[4]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_8 input132 (.A(ref_start_addr[5]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(ref_start_addr[6]),
    .X(net133));
 sky130_fd_sc_hd__buf_8 input134 (.A(ref_start_addr[7]),
    .X(net134));
 sky130_fd_sc_hd__dlymetal6s2s_1 input135 (.A(ref_start_addr[8]),
    .X(net135));
 sky130_fd_sc_hd__buf_4 input136 (.A(ref_start_addr[9]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 input137 (.A(rst_n),
    .X(net137));
 sky130_fd_sc_hd__buf_4 input138 (.A(start),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 output139 (.A(net139),
    .X(done));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(mem_addr[0]));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net141),
    .X(mem_addr[10]));
 sky130_fd_sc_hd__clkbuf_4 output142 (.A(net142),
    .X(mem_addr[11]));
 sky130_fd_sc_hd__clkbuf_4 output143 (.A(net208),
    .X(mem_addr[12]));
 sky130_fd_sc_hd__clkbuf_4 output144 (.A(net207),
    .X(mem_addr[13]));
 sky130_fd_sc_hd__clkbuf_4 output145 (.A(net145),
    .X(mem_addr[14]));
 sky130_fd_sc_hd__clkbuf_4 output146 (.A(net206),
    .X(mem_addr[15]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(mem_addr[16]));
 sky130_fd_sc_hd__clkbuf_4 output148 (.A(net204),
    .X(mem_addr[17]));
 sky130_fd_sc_hd__clkbuf_4 output149 (.A(net149),
    .X(mem_addr[18]));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net150),
    .X(mem_addr[19]));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net151),
    .X(mem_addr[1]));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net201),
    .X(mem_addr[20]));
 sky130_fd_sc_hd__clkbuf_4 output153 (.A(net153),
    .X(mem_addr[21]));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net154),
    .X(mem_addr[22]));
 sky130_fd_sc_hd__clkbuf_4 output155 (.A(net155),
    .X(mem_addr[23]));
 sky130_fd_sc_hd__clkbuf_4 output156 (.A(net156),
    .X(mem_addr[24]));
 sky130_fd_sc_hd__clkbuf_4 output157 (.A(net200),
    .X(mem_addr[25]));
 sky130_fd_sc_hd__clkbuf_4 output158 (.A(net158),
    .X(mem_addr[26]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(mem_addr[27]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(mem_addr[28]));
 sky130_fd_sc_hd__clkbuf_4 output161 (.A(net161),
    .X(mem_addr[29]));
 sky130_fd_sc_hd__clkbuf_4 output162 (.A(net162),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__buf_6 output163 (.A(net163),
    .X(mem_addr[30]));
 sky130_fd_sc_hd__buf_6 output164 (.A(net164),
    .X(mem_addr[31]));
 sky130_fd_sc_hd__clkbuf_4 output165 (.A(net165),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__clkbuf_4 output166 (.A(net166),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__clkbuf_4 output167 (.A(net210),
    .X(mem_addr[5]));
 sky130_fd_sc_hd__clkbuf_4 output168 (.A(net168),
    .X(mem_addr[6]));
 sky130_fd_sc_hd__clkbuf_4 output169 (.A(net169),
    .X(mem_addr[7]));
 sky130_fd_sc_hd__clkbuf_4 output170 (.A(net170),
    .X(mem_addr[8]));
 sky130_fd_sc_hd__clkbuf_4 output171 (.A(net171),
    .X(mem_addr[9]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(mv_x[0]));
 sky130_fd_sc_hd__clkbuf_4 output173 (.A(net173),
    .X(mv_x[1]));
 sky130_fd_sc_hd__clkbuf_4 output174 (.A(net174),
    .X(mv_x[2]));
 sky130_fd_sc_hd__clkbuf_4 output175 (.A(net175),
    .X(mv_x[3]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(mv_x[4]));
 sky130_fd_sc_hd__clkbuf_4 output177 (.A(net177),
    .X(mv_x[5]));
 sky130_fd_sc_hd__clkbuf_4 output178 (.A(net178),
    .X(mv_y[0]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(mv_y[1]));
 sky130_fd_sc_hd__clkbuf_4 output180 (.A(net180),
    .X(mv_y[2]));
 sky130_fd_sc_hd__clkbuf_4 output181 (.A(net181),
    .X(mv_y[3]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(mv_y[4]));
 sky130_fd_sc_hd__clkbuf_4 output183 (.A(net183),
    .X(mv_y[5]));
 sky130_fd_sc_hd__clkbuf_4 output184 (.A(net184),
    .X(sad[0]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(sad[10]));
 sky130_fd_sc_hd__clkbuf_4 output186 (.A(net186),
    .X(sad[11]));
 sky130_fd_sc_hd__clkbuf_4 output187 (.A(net187),
    .X(sad[12]));
 sky130_fd_sc_hd__clkbuf_4 output188 (.A(net188),
    .X(sad[13]));
 sky130_fd_sc_hd__clkbuf_4 output189 (.A(net189),
    .X(sad[14]));
 sky130_fd_sc_hd__clkbuf_4 output190 (.A(net190),
    .X(sad[15]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(sad[1]));
 sky130_fd_sc_hd__clkbuf_4 output192 (.A(net192),
    .X(sad[2]));
 sky130_fd_sc_hd__clkbuf_4 output193 (.A(net193),
    .X(sad[3]));
 sky130_fd_sc_hd__clkbuf_4 output194 (.A(net194),
    .X(sad[4]));
 sky130_fd_sc_hd__clkbuf_4 output195 (.A(net195),
    .X(sad[5]));
 sky130_fd_sc_hd__clkbuf_4 output196 (.A(net196),
    .X(sad[6]));
 sky130_fd_sc_hd__clkbuf_4 output197 (.A(net197),
    .X(sad[7]));
 sky130_fd_sc_hd__clkbuf_4 output198 (.A(net198),
    .X(sad[8]));
 sky130_fd_sc_hd__clkbuf_4 output199 (.A(net199),
    .X(sad[9]));
 sky130_fd_sc_hd__buf_6 wire200 (.A(net157),
    .X(net200));
 sky130_fd_sc_hd__buf_4 wire201 (.A(net152),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 max_cap202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 max_cap203 (.A(_05705_),
    .X(net203));
 sky130_fd_sc_hd__buf_6 wire204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_4 wire205 (.A(net148),
    .X(net205));
 sky130_fd_sc_hd__buf_4 wire206 (.A(net146),
    .X(net206));
 sky130_fd_sc_hd__buf_6 wire207 (.A(net144),
    .X(net207));
 sky130_fd_sc_hd__buf_6 wire208 (.A(net143),
    .X(net208));
 sky130_fd_sc_hd__buf_1 max_cap209 (.A(_05361_),
    .X(net209));
 sky130_fd_sc_hd__buf_4 wire210 (.A(net167),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 wire211 (.A(net2000),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 max_cap212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 wire213 (.A(_04554_),
    .X(net213));
 sky130_fd_sc_hd__buf_6 load_slew214 (.A(_03807_),
    .X(net214));
 sky130_fd_sc_hd__buf_6 load_slew215 (.A(_09123_),
    .X(net215));
 sky130_fd_sc_hd__buf_6 max_cap216 (.A(_08980_),
    .X(net216));
 sky130_fd_sc_hd__buf_4 wire217 (.A(_05885_),
    .X(net217));
 sky130_fd_sc_hd__buf_6 max_cap218 (.A(_02527_),
    .X(net218));
 sky130_fd_sc_hd__buf_1 max_cap219 (.A(net2001),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_8 max_cap220 (.A(_06196_),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_8 max_cap221 (.A(_06176_),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 max_cap222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 max_cap223 (.A(_06078_),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 wire224 (.A(net2003),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 max_cap225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 max_cap226 (.A(_06004_),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 wire227 (.A(net2005),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 max_cap228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 wire229 (.A(net231),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 max_cap230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 max_cap231 (.A(_05992_),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 wire232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 max_cap233 (.A(net235),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 max_cap234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 wire235 (.A(net2006),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 max_cap236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 max_cap237 (.A(net238),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 max_cap238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 max_cap239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 max_cap240 (.A(net241),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 wire241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 wire242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 wire243 (.A(_05969_),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 wire244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 max_cap245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 max_cap246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 wire247 (.A(net249),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 max_cap248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 wire249 (.A(_05932_),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_2 wire250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 max_cap251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_2 max_cap252 (.A(_05926_),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_8 max_cap253 (.A(_05913_),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 max_cap254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 max_cap255 (.A(net259),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_2 max_cap256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_2 max_cap257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 max_cap258 (.A(net2007),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 max_cap259 (.A(_05894_),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_2 wire260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_2 wire261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 wire262 (.A(net265),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 max_cap263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_2 max_cap264 (.A(net2008),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 max_cap265 (.A(net2008),
    .X(net265));
 sky130_fd_sc_hd__buf_4 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__buf_2 fanout267 (.A(net280),
    .X(net267));
 sky130_fd_sc_hd__buf_4 fanout268 (.A(net271),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_4 fanout269 (.A(net271),
    .X(net269));
 sky130_fd_sc_hd__buf_4 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(net280),
    .X(net271));
 sky130_fd_sc_hd__buf_4 fanout272 (.A(net275),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 fanout273 (.A(net275),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 fanout275 (.A(net279),
    .X(net275));
 sky130_fd_sc_hd__buf_4 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_4 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 fanout278 (.A(net280),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_8 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__buf_8 fanout280 (.A(net137),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_227_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_232_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_233_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_252_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_253_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_257_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_258_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_259_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_261_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_262_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_264_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_265_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_268_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_269_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_270_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_271_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_272_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_273_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_274_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_275_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_276_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_276_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_277_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_278_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_279_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_280_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_281_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_282_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_283_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_284_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_285_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_285_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_286_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_286_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_287_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_287_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_288_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_288_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_289_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_289_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_290_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_290_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_291_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_291_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_292_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_292_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_293_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_293_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_294_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_294_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_295_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_295_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_296_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_296_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_297_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_297_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_298_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_298_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_299_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_299_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_300_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_300_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_301_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_301_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_302_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_302_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_303_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_303_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_304_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_304_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_305_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_305_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_306_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_306_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_307_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_307_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_308_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_308_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_309_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_309_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_310_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_310_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_311_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_311_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_312_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_312_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_313_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_313_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_314_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_314_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_315_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_315_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_316_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_316_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_317_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_317_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_318_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_318_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_319_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_319_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_320_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_320_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_321_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_321_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_322_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_322_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_323_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_323_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_324_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_324_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_325_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_325_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_326_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_326_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_327_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_327_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_328_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_328_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_329_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_329_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_330_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_330_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_331_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_331_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_332_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_332_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_333_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_333_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_334_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_334_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_335_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_335_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_336_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_336_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_337_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_337_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_338_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_338_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_339_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_339_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_340_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_340_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_341_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_341_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_342_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_342_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_343_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_343_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_344_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_344_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_345_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_345_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_346_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_346_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_347_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_347_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_348_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_348_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_349_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_349_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_350_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_350_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_351_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_351_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_352_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_352_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_353_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_353_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_354_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_354_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_355_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_355_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_356_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_356_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_357_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_357_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_358_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_358_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_359_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_359_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_360_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_360_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_361_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_361_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_362_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_362_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_363_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_363_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_364_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_364_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_365_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_365_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_366_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_366_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_367_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_367_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_368_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_368_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_369_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_369_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_370_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_370_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_371_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_371_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_372_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_372_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_373_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_373_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_374_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_374_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_375_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_375_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_376_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_376_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_377_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_377_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_378_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_378_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_379_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_379_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_380_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_380_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_381_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_381_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_382_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_382_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_383_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_383_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_384_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_384_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_385_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_385_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_386_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_386_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_387_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_387_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_388_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_388_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_389_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_389_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_390_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_390_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_391_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_391_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_392_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_392_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_393_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_393_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_394_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_394_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_2__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_3__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_4__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_5__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_6__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_7__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_8__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_9__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_10__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_11__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_12__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_13__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_14__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_15__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_15__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_16__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_17__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_18__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_19__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_20__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_21__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_22__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_22__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_23__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_24__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_25__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_26__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_27__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_28__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_29__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_30__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_31__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 rebuffer1 (.A(_05233_),
    .X(net281));
 sky130_fd_sc_hd__buf_1 rebuffer2 (.A(_04795_),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 rebuffer3 (.A(_04934_),
    .X(net283));
 sky130_fd_sc_hd__buf_2 split4 (.A(_04781_),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(_04741_),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 rebuffer6 (.A(net2002),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(_05116_),
    .X(net287));
 sky130_fd_sc_hd__buf_1 rebuffer8 (.A(_04835_),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_1 rebuffer9 (.A(net288),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 rebuffer10 (.A(_04794_),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\best_point_idx[2] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_04446_),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\current_accum_sad[5] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\current_accum_sad[4] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\current_accum_sad[3] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\current_accum_sad[15] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\pixel_cnt[8] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\current_accum_sad[6] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\current_accum_sad[14] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\current_accum_sad[0] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\current_accum_sad[1] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\current_accum_sad[13] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\current_accum_sad[12] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\current_accum_sad[7] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\current_accum_sad[2] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\cand_y[4] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\current_accum_sad[9] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\current_accum_sad[10] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\point_cnt[3] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\state[5] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\cur_mb_mem[89][3] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\cur_mb_mem[188][0] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\cur_mb_mem[153][2] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\cur_mb_mem[170][7] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\cur_mb_mem[86][3] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\cur_mb_mem[108][1] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\cur_mb_mem[93][0] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\cur_mb_mem[111][2] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\cur_mb_mem[188][5] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\cur_mb_mem[57][0] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\cur_mb_mem[170][3] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\cur_mb_mem[86][5] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\cur_mb_mem[188][6] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\cur_mb_mem[174][5] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\cur_mb_mem[165][2] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\cur_mb_mem[183][5] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\cur_mb_mem[101][5] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\cur_mb_mem[105][3] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\cur_mb_mem[103][1] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\cur_mb_mem[109][4] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\cur_mb_mem[58][1] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\cur_mb_mem[93][4] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\cur_mb_mem[229][7] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\cur_mb_mem[111][3] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\cur_mb_mem[171][4] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\cur_mb_mem[89][1] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\cur_mb_mem[252][5] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\cur_mb_mem[252][2] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\cur_mb_mem[155][1] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\cur_mb_mem[179][3] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\cur_mb_mem[117][3] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\cur_mb_mem[172][3] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\cur_mb_mem[60][3] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\cur_mb_mem[109][2] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\cur_mb_mem[181][1] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\cur_mb_mem[89][0] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\cur_mb_mem[87][3] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\cur_mb_mem[54][1] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\cur_mb_mem[105][4] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\cur_mb_mem[147][1] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\cur_mb_mem[103][2] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\cur_mb_mem[165][1] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\cur_mb_mem[188][7] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\cur_mb_mem[93][3] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\cur_mb_mem[174][2] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\cur_mb_mem[92][7] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\cur_mb_mem[106][4] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\cur_mb_mem[7][0] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\cur_mb_mem[126][1] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\cur_mb_mem[87][4] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\cur_mb_mem[174][1] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\cur_mb_mem[93][6] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\cur_mb_mem[163][1] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\cur_mb_mem[86][0] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\cur_mb_mem[254][2] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\cur_mb_mem[115][5] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\cur_mb_mem[237][4] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\cur_mb_mem[7][5] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\cur_mb_mem[90][0] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\cur_mb_mem[187][4] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\cur_mb_mem[173][5] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\cur_mb_mem[154][2] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\cur_mb_mem[87][1] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\cur_mb_mem[99][5] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\cur_mb_mem[179][4] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\cur_mb_mem[90][5] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\cur_mb_mem[59][1] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\cur_mb_mem[92][6] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\cur_mb_mem[111][0] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\cur_mb_mem[175][5] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\cur_mb_mem[90][7] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\cur_mb_mem[169][5] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\cur_mb_mem[171][0] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\cur_mb_mem[252][1] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\cur_mb_mem[57][1] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\cur_mb_mem[117][0] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\cur_mb_mem[125][4] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\cur_mb_mem[102][4] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\state[2] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\cur_mb_mem[7][2] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\cur_mb_mem[173][4] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\cur_mb_mem[93][2] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\cur_mb_mem[57][4] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\cur_mb_mem[172][1] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\cur_mb_mem[179][0] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\cur_mb_mem[193][3] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\cur_mb_mem[63][2] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\best_point_idx[3] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\cur_mb_mem[138][1] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\cur_mb_mem[188][4] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\cur_mb_mem[158][3] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\cur_mb_mem[109][3] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\cur_mb_mem[173][0] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\cur_mb_mem[72][3] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\cur_mb_mem[249][3] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\cur_mb_mem[171][2] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\cur_mb_mem[57][3] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\cur_mb_mem[60][2] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\cur_mb_mem[165][5] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\cur_mb_mem[7][4] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\cur_mb_mem[63][3] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\cur_mb_mem[187][3] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\cur_mb_mem[183][3] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\cur_mb_mem[115][4] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\cur_mb_mem[170][5] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\cur_mb_mem[58][0] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\cur_mb_mem[165][0] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\cur_mb_mem[183][0] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\cur_mb_mem[102][5] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\cur_mb_mem[251][4] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\cur_mb_mem[167][3] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\cur_mb_mem[119][0] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\cur_mb_mem[55][1] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\cur_mb_mem[157][1] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\cur_mb_mem[87][2] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\cur_mb_mem[123][1] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\cur_mb_mem[94][3] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\cur_mb_mem[158][0] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\cur_mb_mem[58][5] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\cur_mb_mem[186][5] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\cur_mb_mem[182][5] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\cur_mb_mem[254][3] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\cur_mb_mem[249][0] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\cur_mb_mem[93][1] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\cur_mb_mem[119][2] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\cur_mb_mem[174][4] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\cur_mb_mem[230][7] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\cur_mb_mem[63][0] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\cur_mb_mem[107][2] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\cur_mb_mem[121][2] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\cur_mb_mem[153][3] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\cur_mb_mem[63][5] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\cur_mb_mem[172][4] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\cur_mb_mem[115][7] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\cur_mb_mem[147][6] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\cur_mb_mem[55][2] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\cur_mb_mem[170][2] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\cur_mb_mem[169][2] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\cur_mb_mem[9][6] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\cur_mb_mem[153][0] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\cur_mb_mem[146][1] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\cur_mb_mem[99][3] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\cur_mb_mem[7][3] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\cur_mb_mem[90][3] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\cur_mb_mem[101][4] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\cur_mb_mem[109][1] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\cur_mb_mem[99][4] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\cur_mb_mem[154][3] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\cur_mb_mem[86][1] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\cur_mb_mem[171][3] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\cur_mb_mem[58][3] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\cur_mb_mem[107][1] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\cur_mb_mem[53][1] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\cur_mb_mem[106][0] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\cur_mb_mem[89][4] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\cur_mb_mem[92][5] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\cur_mb_mem[183][6] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\cur_mb_mem[171][7] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\cur_mb_mem[170][0] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\cur_mb_mem[252][4] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\cur_mb_mem[60][4] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\cur_mb_mem[163][5] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\cur_mb_mem[115][1] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\cur_mb_mem[187][5] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\cur_mb_mem[93][5] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\cur_mb_mem[187][6] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\cur_mb_mem[173][2] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\cur_mb_mem[76][3] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\cur_mb_mem[103][0] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\cur_mb_mem[115][3] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\cur_mb_mem[179][2] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\cur_mb_mem[106][2] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\cur_mb_mem[64][1] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\cur_mb_mem[163][0] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\cur_mb_mem[167][1] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\cur_mb_mem[102][3] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\cur_mb_mem[76][4] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\cur_mb_mem[91][5] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\cur_mb_mem[92][4] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\cur_mb_mem[95][4] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\cur_mb_mem[92][0] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\cur_mb_mem[186][4] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\cur_mb_mem[90][2] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\cur_mb_mem[92][2] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\cur_mb_mem[49][0] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\cur_mb_mem[183][2] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\cur_mb_mem[92][3] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\cur_mb_mem[194][0] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\cur_mb_mem[106][3] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\cur_mb_mem[173][1] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\cur_mb_mem[71][2] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\cur_mb_mem[149][5] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\cur_mb_mem[169][4] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\cur_mb_mem[48][0] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\cur_mb_mem[172][5] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\cur_mb_mem[7][1] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\cur_mb_mem[94][0] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\cur_mb_mem[171][5] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\cur_mb_mem[167][2] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\cur_mb_mem[149][3] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\cur_mb_mem[33][3] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\cur_mb_mem[208][2] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\cur_mb_mem[102][0] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\cur_mb_mem[185][5] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\cur_mb_mem[105][5] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\cur_mb_mem[188][1] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\cur_mb_mem[89][5] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\cur_mb_mem[62][2] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\cur_mb_mem[181][0] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\cur_mb_mem[137][1] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\cur_mb_mem[186][1] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\cur_mb_mem[58][4] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\cur_mb_mem[181][4] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\cur_mb_mem[59][2] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\cur_mb_mem[173][3] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\cur_mb_mem[229][4] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\cur_mb_mem[99][0] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\cur_mb_mem[99][2] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\cur_mb_mem[5][4] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\cur_mb_mem[54][5] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\cur_mb_mem[80][0] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\cur_mb_mem[105][0] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\cur_mb_mem[183][1] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\cur_mb_mem[181][3] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\cur_mb_mem[147][0] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\cur_mb_mem[196][4] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\cur_mb_mem[172][0] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\cur_mb_mem[251][0] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\cur_mb_mem[175][1] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\cur_mb_mem[179][5] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\cur_mb_mem[94][1] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\cur_mb_mem[50][1] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\cur_mb_mem[119][1] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\cur_mb_mem[176][5] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\cur_mb_mem[123][2] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\cur_mb_mem[39][1] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\cur_mb_mem[160][5] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\cur_mb_mem[107][3] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\cur_mb_mem[125][2] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\cur_mb_mem[163][4] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\cur_mb_mem[54][7] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\cur_mb_mem[149][4] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\cur_mb_mem[94][2] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\cur_mb_mem[87][5] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\cur_mb_mem[160][7] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\cur_mb_mem[167][0] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\cur_mb_mem[91][4] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\cur_mb_mem[94][4] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\cur_mb_mem[212][3] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\cur_mb_mem[59][3] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\cur_mb_mem[59][0] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\cur_mb_mem[136][0] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\cur_mb_mem[62][5] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\cur_mb_mem[182][4] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\best_cand_x[6] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\cur_mb_mem[123][0] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\cur_mb_mem[83][7] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\cur_mb_mem[137][0] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\cur_mb_mem[210][3] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\cur_mb_mem[145][3] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\cur_mb_mem[163][2] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\cur_mb_mem[86][4] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\cur_mb_mem[169][1] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\cur_mb_mem[106][1] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\cur_mb_mem[196][1] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\cur_mb_mem[43][0] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\cur_mb_mem[60][0] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\cur_mb_mem[87][0] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\cur_mb_mem[16][3] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\cur_mb_mem[107][4] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\cur_mb_mem[148][5] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\cur_mb_mem[82][0] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\cur_mb_mem[249][5] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\cur_mb_mem[150][0] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\cur_mb_mem[92][1] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\cur_mb_mem[222][1] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\cur_mb_mem[99][1] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\cur_mb_mem[85][7] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\cur_mb_mem[254][0] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\cur_mb_mem[121][0] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\cur_mb_mem[23][0] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\cur_mb_mem[168][0] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\cur_mb_mem[134][4] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\cur_mb_mem[75][4] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\cur_mb_mem[136][1] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\cur_mb_mem[137][3] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\cur_mb_mem[13][1] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\cur_mb_mem[249][2] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\best_point_idx[1] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\cur_mb_mem[59][6] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\cur_mb_mem[37][4] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\cur_mb_mem[209][3] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\cur_mb_mem[171][1] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\cur_mb_mem[186][0] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\cur_mb_mem[123][3] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\cur_mb_mem[230][2] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\cur_mb_mem[130][0] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\cur_mb_mem[139][3] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\cur_mb_mem[252][0] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\cur_mb_mem[60][1] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\cur_mb_mem[251][3] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\cur_mb_mem[27][3] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\cur_mb_mem[82][5] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\cur_mb_mem[18][1] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\cur_mb_mem[230][4] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\cur_mb_mem[76][2] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\cur_mb_mem[76][0] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\cur_mb_mem[48][5] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\cur_mb_mem[169][3] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\cur_mb_mem[16][1] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\cur_mb_mem[162][1] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\cur_mb_mem[91][7] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\current_accum_sad[11] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\cur_mb_mem[55][6] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\cur_mb_mem[54][4] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\cur_mb_mem[34][3] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\cur_mb_mem[139][0] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\cur_mb_mem[18][5] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\cur_mb_mem[181][2] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\cur_mb_mem[105][1] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\cur_mb_mem[94][5] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\cur_mb_mem[142][4] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\cur_mb_mem[149][1] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\cur_mb_mem[49][4] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\cur_mb_mem[210][0] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\cur_mb_mem[192][7] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\cur_mb_mem[160][4] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\cur_mb_mem[109][0] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\cur_mb_mem[13][7] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\cur_mb_mem[236][5] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\cur_mb_mem[220][0] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\cur_mb_mem[57][5] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\cur_mb_mem[83][6] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\cur_mb_mem[107][5] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\cur_mb_mem[88][5] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\cur_mb_mem[148][1] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\cur_mb_mem[121][3] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\cur_mb_mem[62][0] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\cur_mb_mem[49][1] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\cur_mb_mem[102][2] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\cur_mb_mem[183][4] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\cur_mb_mem[247][4] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\cur_mb_mem[81][0] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\cur_mb_mem[48][4] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\cur_mb_mem[77][4] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\cur_mb_mem[59][4] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\cur_mb_mem[17][1] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\cur_mb_mem[122][3] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\cur_mb_mem[124][6] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\cur_mb_mem[165][4] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\cur_mb_mem[181][5] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\cur_mb_mem[134][5] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\cur_mb_mem[40][0] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\cur_mb_mem[136][3] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\cur_mb_mem[170][4] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\cur_mb_mem[144][4] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\cur_mb_mem[200][0] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\cur_mb_mem[210][5] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\cur_mb_mem[63][4] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\cur_mb_mem[1][3] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\cur_mb_mem[174][3] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\cur_mb_mem[109][5] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\cur_mb_mem[132][1] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\cur_mb_mem[16][5] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\cur_mb_mem[52][1] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\cur_mb_mem[3][0] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\cur_mb_mem[255][6] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\cur_mb_mem[51][3] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\cur_mb_mem[82][2] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\cur_mb_mem[147][3] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\cur_mb_mem[184][3] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\cur_mb_mem[229][1] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\cur_mb_mem[64][3] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\cur_mb_mem[62][3] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\cur_mb_mem[76][5] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\cur_mb_mem[17][0] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\cur_mb_mem[137][5] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\cur_mb_mem[117][2] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\cur_mb_mem[122][7] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\cur_mb_mem[163][3] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\cur_mb_mem[78][0] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\cur_mb_mem[126][3] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\cur_mb_mem[75][5] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\cur_mb_mem[9][4] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\cur_mb_mem[172][2] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\cur_mb_mem[55][0] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\cur_mb_mem[102][7] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\best_cand_y[6] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\cur_mb_mem[255][1] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\cur_mb_mem[185][4] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\cur_mb_mem[36][5] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\cur_mb_mem[240][2] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\cur_mb_mem[220][4] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\cur_mb_mem[43][2] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\cur_mb_mem[68][4] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\cur_mb_mem[237][5] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\cur_mb_mem[56][5] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\cur_mb_mem[84][4] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\cur_mb_mem[140][1] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\cur_mb_mem[171][6] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\cur_mb_mem[48][3] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\cur_mb_mem[47][2] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\cur_mb_mem[49][5] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\cur_mb_mem[54][3] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\cur_mb_mem[43][3] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\cur_mb_mem[9][1] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\cur_mb_mem[159][6] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\cur_mb_mem[35][4] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\cur_mb_mem[194][3] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\cur_mb_mem[21][2] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\cur_mb_mem[196][5] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\cur_mb_mem[196][2] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\cur_mb_mem[69][0] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\cur_mb_mem[133][2] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\cur_mb_mem[255][4] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\cur_mb_mem[142][5] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\best_point_idx[0] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\cur_mb_mem[6][4] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\cur_mb_mem[251][2] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\cur_mb_mem[200][2] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\cur_mb_mem[131][1] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\cur_mb_mem[126][0] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\cur_mb_mem[129][4] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\cur_mb_mem[5][5] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\cur_mb_mem[94][6] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\cur_mb_mem[64][4] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\cur_mb_mem[71][4] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\cur_mb_mem[34][0] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\cur_mb_mem[16][0] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\cur_mb_mem[13][6] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\cur_mb_mem[88][4] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\cur_mb_mem[119][7] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\cur_mb_mem[77][3] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\cur_mb_mem[220][1] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\cur_mb_mem[145][4] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\cur_mb_mem[126][2] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\cur_mb_mem[133][3] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\cur_mb_mem[125][3] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\cur_mb_mem[177][5] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\cur_mb_mem[208][1] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\cur_mb_mem[220][5] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\cur_mb_mem[49][2] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\cur_mb_mem[187][2] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\cur_mb_mem[14][6] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\cur_mb_mem[90][4] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\cur_mb_mem[254][6] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\cur_mb_mem[227][5] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\cur_mb_mem[165][3] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\cur_mb_mem[147][7] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\cur_mb_mem[168][4] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\cur_mb_mem[57][7] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\cur_mb_mem[85][3] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\cur_mb_mem[155][5] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\cur_mb_mem[44][5] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\cur_mb_mem[144][5] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\cur_mb_mem[91][3] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\cur_mb_mem[168][2] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\cur_mb_mem[178][3] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\cur_mb_mem[188][3] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\cur_mb_mem[175][4] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\cur_mb_mem[244][3] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\cur_mb_mem[49][3] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\cur_mb_mem[84][3] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\cur_mb_mem[170][1] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\cur_mb_mem[41][2] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\cur_mb_mem[130][5] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\cur_mb_mem[254][4] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\cur_mb_mem[84][1] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\cur_mb_mem[23][3] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\cur_mb_mem[166][1] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\cur_mb_mem[145][0] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\cur_mb_mem[130][4] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\cur_mb_mem[63][1] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\cur_mb_mem[186][2] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\cur_mb_mem[110][3] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\cur_mb_mem[111][4] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\cur_mb_mem[52][5] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\cur_mb_mem[135][1] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\cur_mb_mem[106][7] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\cur_mb_mem[210][4] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\cur_mb_mem[60][7] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\cur_mb_mem[17][2] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\cur_mb_mem[21][3] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\cur_mb_mem[193][0] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\cur_mb_mem[222][7] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\cur_mb_mem[91][6] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\cur_mb_mem[250][5] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\cur_mb_mem[146][0] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\cur_mb_mem[35][5] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\cur_mb_mem[14][1] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\cur_mb_mem[20][1] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\cur_mb_mem[84][5] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\cur_mb_mem[156][7] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\cur_mb_mem[221][7] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\cur_mb_mem[39][4] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\cur_mb_mem[40][3] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\cur_mb_mem[85][1] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\cur_mb_mem[192][1] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\cur_mb_mem[95][5] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\cur_mb_mem[16][4] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\cur_mb_mem[131][5] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\cur_mb_mem[62][4] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\cur_mb_mem[110][7] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\cur_mb_mem[237][0] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\cur_mb_mem[55][3] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\cur_mb_mem[149][7] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\cur_mb_mem[229][0] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\cur_mb_mem[111][6] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\cur_mb_mem[157][3] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\cur_mb_mem[162][0] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\cur_mb_mem[137][4] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\cur_mb_mem[18][4] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\cur_mb_mem[90][1] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\cur_mb_mem[110][1] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\cur_mb_mem[138][5] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\cur_mb_mem[247][5] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\cur_mb_mem[124][5] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\cur_mb_mem[229][3] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\cur_mb_mem[174][7] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\cur_mb_mem[139][4] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\cur_mb_mem[22][4] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\cur_mb_mem[220][2] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\cur_mb_mem[48][2] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\cur_mb_mem[162][3] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\cur_mb_mem[48][1] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\cur_mb_mem[233][6] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\cur_mb_mem[108][4] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\cur_mb_mem[23][1] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\cur_mb_mem[11][7] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\cur_mb_mem[56][4] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\cur_mb_mem[24][5] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\cur_mb_mem[175][6] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\cur_mb_mem[148][4] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\cur_mb_mem[77][0] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\cur_mb_mem[174][6] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\cur_mb_mem[176][1] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\cur_mb_mem[78][3] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\cur_mb_mem[78][5] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\cur_mb_mem[125][6] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\cur_mb_mem[87][6] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\cur_mb_mem[182][2] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\cur_mb_mem[156][5] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\cur_mb_mem[150][1] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\cur_mb_mem[103][3] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\cur_mb_mem[181][6] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\cur_mb_mem[81][1] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\cur_mb_mem[178][0] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\cur_mb_mem[127][6] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\cur_mb_mem[109][7] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\cur_mb_mem[9][0] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\cur_mb_mem[78][6] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\cur_mb_mem[21][0] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\cur_mb_mem[169][6] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\cur_mb_mem[62][6] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\cur_mb_mem[230][5] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\cur_mb_mem[161][4] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\cur_mb_mem[46][0] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\cur_mb_mem[15][3] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\cur_mb_mem[182][3] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\cur_mb_mem[41][0] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\cur_mb_mem[91][0] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\cur_mb_mem[82][1] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\cur_mb_mem[101][6] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\cur_mb_mem[229][2] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\cur_mb_mem[182][0] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\cur_mb_mem[127][7] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\cur_mb_mem[88][3] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\cur_mb_mem[187][7] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\cur_mb_mem[68][5] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\cur_mb_mem[166][7] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\cur_mb_mem[2][3] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\cur_mb_mem[37][5] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\cur_mb_mem[95][6] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\cur_mb_mem[86][6] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\cur_mb_mem[110][4] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\cur_mb_mem[101][0] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\cur_mb_mem[8][7] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\cur_mb_mem[9][7] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\cur_mb_mem[160][0] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\cur_mb_mem[180][5] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\cur_mb_mem[99][6] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\cur_mb_mem[101][7] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\cur_mb_mem[150][7] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\cur_mb_mem[253][6] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\cur_mb_mem[125][5] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\cur_mb_mem[59][5] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\cur_mb_mem[15][0] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\cur_mb_mem[36][4] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\cur_mb_mem[172][7] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\cur_mb_mem[95][2] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\cur_mb_mem[103][5] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\cur_mb_mem[101][2] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\cur_mb_mem[186][7] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\cur_mb_mem[64][0] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\cur_mb_mem[81][5] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\cur_mb_mem[177][1] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\cur_mb_mem[212][2] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\cur_mb_mem[3][3] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\cur_mb_mem[73][1] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\cur_mb_mem[99][7] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\cur_mb_mem[212][1] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\cur_mb_mem[8][4] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\cur_mb_mem[23][2] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\cur_mb_mem[217][4] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\cur_mb_mem[9][3] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\cur_mb_mem[184][4] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\cur_mb_mem[89][2] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\cur_mb_mem[107][6] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\cur_mb_mem[156][1] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\cur_mb_mem[111][5] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\cur_mb_mem[156][4] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\cur_mb_mem[233][4] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\cur_mb_mem[222][2] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\cur_mb_mem[82][4] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\cur_mb_mem[11][0] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\cur_mb_mem[138][4] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\cur_mb_mem[141][4] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\cur_mb_mem[53][2] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\cur_mb_mem[187][1] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\cur_mb_mem[22][5] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\cur_mb_mem[154][7] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\cur_mb_mem[18][2] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\cur_mb_mem[69][1] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\cur_mb_mem[91][2] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\cur_mb_mem[14][3] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\cur_mb_mem[129][5] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\cur_mb_mem[89][7] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\cur_mb_mem[58][2] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\cur_mb_mem[75][2] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\cur_mb_mem[167][6] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\cur_mb_mem[192][2] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\cur_mb_mem[159][4] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\cur_mb_mem[61][6] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\cur_mb_mem[183][7] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\cur_mb_mem[101][1] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\cur_mb_mem[253][4] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\cur_mb_mem[44][4] ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\cur_mb_mem[243][4] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\cur_mb_mem[227][7] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\cur_mb_mem[185][7] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\cur_mb_mem[28][5] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\cur_mb_mem[224][0] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\cur_mb_mem[184][5] ),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\cur_mb_mem[77][5] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\cur_mb_mem[56][1] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\cur_mb_mem[130][1] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\cur_mb_mem[249][4] ),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\cur_mb_mem[106][5] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\cur_mb_mem[253][7] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\cur_mb_mem[46][4] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\cur_mb_mem[79][1] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\cur_mb_mem[133][1] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\cur_mb_mem[103][7] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\cur_mb_mem[163][6] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\cur_mb_mem[144][1] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\cur_mb_mem[150][4] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\cur_mb_mem[55][7] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\cur_mb_mem[121][5] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\cur_mb_mem[3][5] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\cur_mb_mem[127][4] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\cur_mb_mem[130][2] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\cur_mb_mem[154][6] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\cur_mb_mem[30][1] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\cur_mb_mem[169][7] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\best_cand_y[0] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\cur_mb_mem[85][5] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\cur_mb_mem[194][4] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\cur_mb_mem[35][0] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\cur_mb_mem[70][2] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\cur_mb_mem[169][0] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\cur_mb_mem[151][1] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\cur_mb_mem[67][1] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\cur_mb_mem[212][5] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\cur_mb_mem[177][4] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\cur_mb_mem[88][2] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\cur_mb_mem[166][2] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\cur_mb_mem[82][7] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\cur_mb_mem[118][3] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\cur_mb_mem[146][2] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\cur_mb_mem[122][2] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\cur_mb_mem[230][6] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\cur_mb_mem[40][2] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\cur_mb_mem[103][4] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\cur_mb_mem[61][5] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\cur_mb_mem[165][6] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\cur_mb_mem[24][4] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\cur_mb_mem[23][5] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\cur_mb_mem[175][2] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\cur_mb_mem[53][7] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\cur_mb_mem[119][3] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\cur_mb_mem[131][4] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\cur_mb_mem[70][3] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\cur_mb_mem[66][6] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\cur_mb_mem[78][4] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\cur_mb_mem[61][7] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\cur_mb_mem[63][6] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\cur_mb_mem[6][1] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\cur_mb_mem[20][6] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\cur_mb_mem[81][3] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\cur_mb_mem[35][3] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\cur_mb_mem[118][6] ),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\cur_mb_mem[53][5] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\cur_mb_mem[158][1] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\cur_mb_mem[157][7] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\cur_mb_mem[179][1] ),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\cur_mb_mem[14][7] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\cur_mb_mem[170][6] ),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\cur_mb_mem[160][3] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\cur_mb_mem[161][5] ),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\cur_mb_mem[58][6] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\cur_mb_mem[143][4] ),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\cur_mb_mem[130][3] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\cur_mb_mem[94][7] ),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\cur_mb_mem[180][4] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\cur_mb_mem[168][1] ),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\cur_mb_mem[147][2] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\cur_mb_mem[6][5] ),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\cur_mb_mem[208][7] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\cur_mb_mem[137][2] ),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\cur_mb_mem[72][7] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\cur_mb_mem[60][5] ),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\cur_mb_mem[208][4] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\cur_mb_mem[157][6] ),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\cur_mb_mem[118][4] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\cur_mb_mem[250][0] ),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\cur_mb_mem[8][3] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\cur_mb_mem[167][7] ),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\cur_mb_mem[51][5] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\cur_mb_mem[51][1] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\cur_mb_mem[219][1] ),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\cur_mb_mem[127][2] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\cur_mb_mem[178][5] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\cur_mb_mem[14][5] ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\cur_mb_mem[34][2] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\cur_mb_mem[192][6] ),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\cur_mb_mem[251][5] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\cur_mb_mem[78][1] ),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\cur_mb_mem[192][5] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\cur_mb_mem[107][0] ),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\cur_mb_mem[58][7] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\cur_mb_mem[105][7] ),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\cur_mb_mem[180][1] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\cur_mb_mem[208][3] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\cur_mb_mem[82][3] ),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\cur_mb_mem[65][3] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\cur_mb_mem[160][1] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\cur_mb_mem[164][7] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\cur_mb_mem[121][1] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\cur_mb_mem[141][5] ),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\cur_mb_mem[65][0] ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\cur_mb_mem[6][2] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\cur_mb_mem[173][6] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\cur_mb_mem[178][1] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\cur_mb_mem[60][6] ),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\cur_mb_mem[52][4] ),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\cur_mb_mem[93][7] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\cur_mb_mem[159][0] ),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\cur_mb_mem[252][3] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\cur_mb_mem[163][7] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\cur_mb_mem[194][7] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\cur_mb_mem[103][6] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\cur_mb_mem[57][6] ),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\cur_mb_mem[182][7] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\cur_mb_mem[250][7] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\cur_mb_mem[166][0] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\cur_mb_mem[179][6] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\cur_mb_mem[86][7] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\cur_mb_mem[21][4] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\cur_mb_mem[9][5] ),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\cur_mb_mem[185][6] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\cur_mb_mem[144][7] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\cur_mb_mem[109][6] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\cur_mb_mem[53][0] ),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\cur_mb_mem[110][2] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\cur_mb_mem[15][6] ),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\cur_mb_mem[132][0] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\cur_mb_mem[161][1] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\cur_mb_mem[209][0] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\cur_mb_mem[254][5] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\cur_mb_mem[23][4] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\cur_mb_mem[70][0] ),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\cur_mb_mem[37][0] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\cur_mb_mem[146][3] ),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\cur_mb_mem[173][7] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\cur_mb_mem[118][5] ),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\cur_mb_mem[182][6] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\cur_mb_mem[140][2] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\cur_mb_mem[64][2] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\cur_mb_mem[39][5] ),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\cur_mb_mem[152][2] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\cur_mb_mem[21][7] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(\cur_mb_mem[127][3] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\cur_mb_mem[76][1] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\cur_mb_mem[251][7] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\cur_mb_mem[211][4] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\cur_mb_mem[69][3] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\cur_mb_mem[75][7] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\cur_mb_mem[221][6] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\cur_mb_mem[152][6] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\cur_mb_mem[145][5] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\cur_mb_mem[227][4] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\cur_mb_mem[162][6] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\cur_mb_mem[255][5] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\cur_mb_mem[186][6] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\cur_mb_mem[149][0] ),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\cur_mb_mem[64][5] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\cur_mb_mem[62][7] ),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\cur_mb_mem[121][4] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\cur_mb_mem[217][3] ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\cur_mb_mem[47][0] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\cur_mb_mem[61][4] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\cur_mb_mem[212][4] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\cur_mb_mem[150][2] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\cur_mb_mem[18][6] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\cur_mb_mem[166][4] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\cur_mb_mem[193][4] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\cur_mb_mem[222][3] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\cur_mb_mem[111][7] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\cur_mb_mem[139][5] ),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\cur_mb_mem[80][3] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\cur_mb_mem[174][0] ),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\cur_mb_mem[102][1] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\cur_mb_mem[175][7] ),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\cur_mb_mem[8][1] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\cur_mb_mem[141][3] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\cur_mb_mem[41][7] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\cur_mb_mem[159][7] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\cur_mb_mem[127][0] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\cur_mb_mem[61][2] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\cur_mb_mem[161][3] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\cur_mb_mem[95][0] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\cur_mb_mem[14][0] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\cur_mb_mem[210][2] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\cur_mb_mem[36][7] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\cur_mb_mem[238][4] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\cur_mb_mem[50][3] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\cur_mb_mem[194][5] ),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\cur_mb_mem[176][4] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\cur_mb_mem[248][7] ),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\cur_mb_mem[42][2] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\cur_mb_mem[236][4] ),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\cur_mb_mem[12][7] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\cur_mb_mem[33][7] ),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\cur_mb_mem[118][1] ),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\cur_mb_mem[43][5] ),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\cur_mb_mem[144][6] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\cur_mb_mem[55][4] ),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\cur_mb_mem[138][7] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\cur_mb_mem[164][5] ),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\cur_mb_mem[8][5] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\cur_mb_mem[193][6] ),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(\cur_mb_mem[253][1] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\cur_mb_mem[19][6] ),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(\cur_mb_mem[42][5] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\cur_mb_mem[142][0] ),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\cur_mb_mem[16][6] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\cur_mb_mem[166][6] ),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\cur_mb_mem[41][5] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\cur_mb_mem[80][2] ),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(\cur_mb_mem[194][2] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\cur_mb_mem[20][0] ),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\cur_mb_mem[34][4] ),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\cur_mb_mem[164][4] ),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(\cur_mb_mem[129][0] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\cur_mb_mem[36][2] ),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\cur_mb_mem[209][2] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\cur_mb_mem[176][7] ),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\cur_mb_mem[63][7] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\cur_mb_mem[130][6] ),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\cur_mb_mem[166][5] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\cur_mb_mem[254][7] ),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(\cur_mb_mem[196][0] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\cur_mb_mem[146][4] ),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\cur_mb_mem[210][6] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\cur_mb_mem[172][6] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(\cur_mb_mem[167][4] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\cur_mb_mem[19][4] ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\cur_mb_mem[36][3] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\cur_mb_mem[155][4] ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\cur_mb_mem[52][2] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\cur_mb_mem[40][1] ),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(\cur_mb_mem[124][2] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\cur_mb_mem[34][6] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\cur_mb_mem[161][7] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\cur_mb_mem[184][7] ),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(\cur_mb_mem[46][1] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\cur_mb_mem[119][6] ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(\cur_mb_mem[10][6] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\cur_mb_mem[48][7] ),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(\cur_mb_mem[145][2] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\cur_mb_mem[162][2] ),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\cur_mb_mem[12][1] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\cur_mb_mem[20][4] ),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(\cur_mb_mem[162][7] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\cur_mb_mem[210][1] ),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\cur_mb_mem[82][6] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\cur_mb_mem[108][5] ),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\cur_mb_mem[3][4] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\cur_mb_mem[35][7] ),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\cur_mb_mem[50][7] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\cur_mb_mem[53][3] ),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\cur_mb_mem[12][5] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\cur_mb_mem[156][6] ),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(\cur_mb_mem[138][3] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\cur_mb_mem[13][5] ),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\cur_mb_mem[0][2] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\cur_mb_mem[145][6] ),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\cur_mb_mem[123][7] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\cur_mb_mem[148][7] ),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\cur_mb_mem[66][5] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\cur_mb_mem[37][7] ),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\cur_mb_mem[143][6] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\cur_mb_mem[253][5] ),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\cur_mb_mem[34][7] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\cur_mb_mem[20][2] ),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\cur_mb_mem[10][2] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\cur_mb_mem[18][0] ),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\cur_mb_mem[72][4] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\cur_mb_mem[42][3] ),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\cur_mb_mem[159][2] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\cur_mb_mem[187][0] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(\cur_mb_mem[44][0] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\cur_mb_mem[38][1] ),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\cur_mb_mem[5][7] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\cur_mb_mem[175][0] ),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\cur_mb_mem[176][2] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\cur_mb_mem[155][2] ),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\cur_mb_mem[164][6] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\cur_mb_mem[137][7] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\cur_mb_mem[85][6] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\cur_mb_mem[139][2] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\cur_mb_mem[141][6] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\cur_mb_mem[66][7] ),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\cur_mb_mem[12][4] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\cur_mb_mem[132][2] ),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\cur_mb_mem[22][7] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\cur_mb_mem[44][1] ),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\cur_mb_mem[210][7] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\cur_mb_mem[86][2] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\cur_mb_mem[255][7] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\cur_mb_mem[226][0] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\cur_mb_mem[178][6] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\cur_mb_mem[151][4] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\cur_mb_mem[75][1] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\cur_mb_mem[7][6] ),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(\cur_mb_mem[151][7] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\cur_mb_mem[139][1] ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(\cur_mb_mem[56][0] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\cur_mb_mem[124][4] ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(\cur_mb_mem[9][2] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\cur_mb_mem[122][0] ),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(\cur_mb_mem[150][5] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\cur_mb_mem[51][6] ),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(\cur_mb_mem[178][4] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\cur_mb_mem[194][1] ),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(\cur_mb_mem[55][5] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\cur_mb_mem[18][7] ),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(\cur_mb_mem[141][7] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\cur_mb_mem[124][0] ),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(\cur_mb_mem[250][2] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\cur_mb_mem[47][3] ),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(\cur_mb_mem[145][7] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\cur_mb_mem[180][6] ),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(\cur_mb_mem[21][6] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\cur_mb_mem[19][7] ),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(\cur_mb_mem[152][5] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\cur_mb_mem[44][3] ),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(\cur_mb_mem[19][2] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\cur_mb_mem[193][2] ),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(\cur_mb_mem[66][3] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\cur_mb_mem[71][5] ),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(\cur_mb_mem[52][3] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\cur_mb_mem[34][5] ),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(\cur_mb_mem[200][4] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\cur_mb_mem[128][0] ),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(\cur_mb_mem[38][4] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\cur_mb_mem[127][1] ),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(\cur_mb_mem[84][7] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\cur_mb_mem[138][0] ),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(\cur_mb_mem[22][1] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\cur_mb_mem[11][5] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(\cur_mb_mem[179][7] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\cur_mb_mem[118][7] ),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(\cur_mb_mem[51][4] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\cur_mb_mem[49][6] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(\cur_mb_mem[231][5] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\cur_mb_mem[225][1] ),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(\cur_mb_mem[51][0] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\cur_mb_mem[139][7] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(\cur_mb_mem[196][3] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\cur_mb_mem[148][6] ),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(\cur_mb_mem[132][3] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\cur_mb_mem[226][2] ),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(\cur_mb_mem[5][6] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\cur_mb_mem[15][1] ),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(\cur_mb_mem[140][5] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\cur_mb_mem[252][6] ),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(\cur_mb_mem[46][5] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\cur_mb_mem[42][6] ),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(\cur_mb_mem[61][1] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\cur_mb_mem[8][0] ),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(\cur_mb_mem[212][7] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\cur_mb_mem[152][4] ),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(\cur_mb_mem[43][6] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\cur_mb_mem[39][3] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(\cur_mb_mem[249][7] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\cur_mb_mem[81][6] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(\cur_mb_mem[36][0] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\cur_mb_mem[175][3] ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(\cur_mb_mem[193][7] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\cur_mb_mem[208][6] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(\cur_mb_mem[136][2] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\cur_mb_mem[143][1] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(\cur_mb_mem[142][1] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\cur_mb_mem[101][3] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(\cur_mb_mem[251][1] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\cur_mb_mem[150][3] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(\cur_mb_mem[89][6] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\cur_mb_mem[49][7] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(\cur_mb_mem[208][0] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\cur_mb_mem[34][1] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(\cur_mb_mem[72][5] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\cur_mb_mem[141][0] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(\cur_mb_mem[22][6] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\cur_mb_mem[15][2] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(\cur_mb_mem[128][5] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\cur_mb_mem[14][4] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(\cur_mb_mem[168][3] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\cur_mb_mem[90][6] ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(\cur_mb_mem[95][1] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\cur_mb_mem[152][0] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(\cur_mb_mem[142][2] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\cur_mb_mem[2][0] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(\cur_mb_mem[167][5] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\cur_mb_mem[110][6] ),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(\cur_mb_mem[226][3] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\cur_mb_mem[79][6] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(\cur_mb_mem[6][7] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\cur_mb_mem[4][4] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(\cur_mb_mem[21][1] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\cur_mb_mem[176][3] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(\cur_mb_mem[56][2] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\cur_mb_mem[139][6] ),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(\cur_mb_mem[138][2] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\cur_mb_mem[13][4] ),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(\cur_mb_mem[152][1] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\cur_mb_mem[228][7] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(\cur_mb_mem[88][7] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\cur_mb_mem[10][7] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(\cur_mb_mem[39][0] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\cur_mb_mem[166][3] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(\cur_mb_mem[75][0] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\cur_mb_mem[6][6] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(\cur_mb_mem[217][5] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\cur_mb_mem[135][5] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(\cur_mb_mem[180][3] ),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\cur_mb_mem[133][0] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(\cur_mb_mem[72][6] ),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\cur_mb_mem[66][4] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(\cur_mb_mem[11][3] ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\cur_mb_mem[43][1] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(\cur_mb_mem[141][1] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\cur_mb_mem[3][6] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(\cur_mb_mem[248][6] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\cur_mb_mem[162][5] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(\cur_mb_mem[8][2] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\cur_mb_mem[25][5] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(\cur_mb_mem[66][1] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\cur_mb_mem[19][0] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(\cur_mb_mem[165][7] ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\cur_mb_mem[248][0] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(\cur_mb_mem[77][7] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\cur_mb_mem[95][7] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(\cur_mb_mem[243][5] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\cur_mb_mem[61][3] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(\cur_mb_mem[46][3] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\cur_mb_mem[108][7] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(\cur_mb_mem[194][6] ),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\cur_mb_mem[178][7] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(\cur_mb_mem[135][4] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\cur_mb_mem[62][1] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(\cur_mb_mem[192][3] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\cur_mb_mem[16][2] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(\cur_mb_mem[17][3] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\cur_mb_mem[19][5] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(\cur_mb_mem[11][2] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\cur_mb_mem[38][5] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(\cur_mb_mem[40][6] ),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\cur_mb_mem[118][0] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(\cur_mb_mem[3][2] ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\cur_mb_mem[158][2] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(\min_sad_reg[8] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\cur_mb_mem[160][2] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(\cur_mb_mem[4][0] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\cur_mb_mem[8][6] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(\cur_mb_mem[142][3] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\cur_mb_mem[95][3] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(\cur_mb_mem[133][6] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\cur_mb_mem[154][5] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(\cur_mb_mem[149][2] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\cur_mb_mem[161][0] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(\cur_mb_mem[17][7] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\cur_mb_mem[78][7] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(\cur_mb_mem[30][0] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\cur_mb_mem[40][4] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(\cur_mb_mem[158][4] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\cur_mb_mem[248][5] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(\cur_mb_mem[37][3] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\cur_mb_mem[48][6] ),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(\cur_mb_mem[143][5] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\cur_mb_mem[116][5] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(\cur_mb_mem[250][3] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\cur_mb_mem[42][4] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(\cur_mb_mem[17][4] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\cur_mb_mem[66][2] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(\cur_mb_mem[15][7] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\cur_mb_mem[200][6] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(\cur_mb_mem[44][6] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(\cur_mb_mem[129][3] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(\cur_mb_mem[145][1] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\cur_mb_mem[10][4] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(\cur_mb_mem[43][4] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\cur_mb_mem[45][2] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(\cur_mb_mem[141][2] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\cur_mb_mem[200][1] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(\cur_mb_mem[220][7] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\cur_mb_mem[106][6] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(\cur_mb_mem[41][4] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(\cur_mb_mem[10][0] ),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(\cur_mb_mem[110][5] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\cur_mb_mem[134][1] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(\cur_mb_mem[64][7] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(\cur_mb_mem[192][0] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(\cur_mb_mem[19][3] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\cur_mb_mem[168][6] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(\cur_mb_mem[11][4] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\cur_mb_mem[146][6] ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(\cur_mb_mem[160][6] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\cur_mb_mem[44][7] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(\cur_mb_mem[132][7] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\cur_mb_mem[154][4] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(\cur_mb_mem[164][2] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\cur_mb_mem[116][4] ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(\cur_mb_mem[46][2] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\cur_mb_mem[161][6] ),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(\cur_mb_mem[31][0] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\cur_mb_mem[28][6] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(\cur_mb_mem[248][4] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\min_sad_reg[4] ),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(\cur_mb_mem[45][0] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\cur_mb_mem[140][4] ),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(\cur_mb_mem[37][1] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\cur_mb_mem[85][2] ),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(\cur_mb_mem[19][1] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\cur_mb_mem[168][7] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(\cur_mb_mem[36][6] ),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\cur_mb_mem[159][3] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(\cur_mb_mem[125][0] ),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\cur_mb_mem[178][2] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(\cur_mb_mem[243][0] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\cur_mb_mem[140][6] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(\cur_mb_mem[200][7] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\cur_mb_mem[185][1] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(\cur_mb_mem[162][4] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\cur_mb_mem[1][5] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(\cur_mb_mem[17][5] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\cur_mb_mem[112][4] ),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(\cur_mb_mem[250][1] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\cur_mb_mem[180][0] ),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(\cur_mb_mem[6][0] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\cur_mb_mem[137][6] ),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(\cur_mb_mem[65][2] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\cur_mb_mem[20][5] ),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(\cur_mb_mem[180][2] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\cur_mb_mem[146][5] ),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(\cur_mb_mem[225][4] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\cur_mb_mem[52][0] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(\cur_mb_mem[38][3] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(\cur_mb_mem[176][0] ),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(\cur_mb_mem[41][3] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\cur_mb_mem[147][4] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(\cur_mb_mem[83][3] ),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\cur_mb_mem[22][3] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(\cur_mb_mem[154][0] ),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\cur_mb_mem[151][5] ),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(\cur_mb_mem[113][5] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\cur_mb_mem[10][5] ),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(\cur_mb_mem[164][3] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\cur_mb_mem[23][7] ),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(\cur_mb_mem[37][6] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\cur_mb_mem[56][3] ),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(\cur_mb_mem[46][6] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\cur_mb_mem[10][1] ),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(\cur_mb_mem[157][0] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\cur_mb_mem[26][0] ),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(\cur_mb_mem[87][7] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\cur_mb_mem[140][7] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(\cur_mb_mem[136][7] ),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\cur_mb_mem[222][0] ),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(\cur_mb_mem[131][6] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\min_sad_reg[3] ),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(\cur_mb_mem[85][4] ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\cur_mb_mem[128][6] ),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(\cur_mb_mem[20][3] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\cur_mb_mem[29][4] ),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(\cur_mb_mem[80][6] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\cur_mb_mem[184][1] ),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(\cur_mb_mem[21][5] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\cur_mb_mem[110][0] ),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(\cur_mb_mem[158][5] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\cur_mb_mem[129][1] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(\cur_mb_mem[211][5] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\cur_mb_mem[225][5] ),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(\cur_mb_mem[6][3] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\cur_mb_mem[238][5] ),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(\cur_mb_mem[75][3] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\cur_mb_mem[143][7] ),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(\cur_mb_mem[250][4] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\cur_mb_mem[71][0] ),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(\cur_mb_mem[16][7] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\cur_mb_mem[25][4] ),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(\cur_mb_mem[77][1] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\cur_mb_mem[164][0] ),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(\cur_mb_mem[22][2] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\cur_mb_mem[42][0] ),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(\cur_mb_mem[38][0] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\cur_mb_mem[76][6] ),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(\cur_mb_mem[47][6] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\cur_mb_mem[32][0] ),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(\cur_mb_mem[24][1] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\cur_mb_mem[242][2] ),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(\cur_mb_mem[43][7] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\cur_mb_mem[227][3] ),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(\cur_mb_mem[248][2] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\cur_mb_mem[2][6] ),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(\cur_mb_mem[52][7] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\cur_mb_mem[35][6] ),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(\cur_mb_mem[196][6] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\cur_mb_mem[128][2] ),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(\cur_mb_mem[108][6] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\cur_mb_mem[3][1] ),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(\cur_mb_mem[220][3] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\cur_mb_mem[193][5] ),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(\cur_mb_mem[67][5] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(\cur_mb_mem[29][5] ),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(\cur_mb_mem[177][6] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(\cur_mb_mem[96][1] ),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(\cur_mb_mem[44][2] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(\cur_mb_mem[38][2] ),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(\cur_mb_mem[78][2] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(\cur_mb_mem[216][2] ),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(\cur_mb_mem[224][5] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\cur_mb_mem[157][5] ),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(\cur_mb_mem[113][2] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(\cur_mb_mem[7][7] ),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(\cur_mb_mem[229][5] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(\cur_mb_mem[67][6] ),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(\cur_mb_mem[27][4] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(\best_cand_y[1] ),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(_00080_),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(\cur_mb_mem[39][6] ),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(\cur_mb_mem[117][5] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(\cur_mb_mem[30][4] ),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(\cur_mb_mem[224][7] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(\cur_mb_mem[40][7] ),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(\cur_mb_mem[2][5] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(\cur_mb_mem[251][6] ),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(\cur_mb_mem[2][2] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(\cur_mb_mem[184][6] ),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(\cur_mb_mem[83][2] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(\min_sad_reg[11] ),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(\cur_mb_mem[161][2] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(\cur_mb_mem[136][5] ),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(\cur_mb_mem[129][2] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(\cur_mb_mem[177][2] ),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(\cur_mb_mem[152][3] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(\cur_mb_mem[81][4] ),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(\cur_mb_mem[2][4] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(\cur_mb_mem[22][0] ),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(\cur_mb_mem[113][4] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(\cur_mb_mem[20][7] ),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(\cur_mb_mem[40][5] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(\cur_mb_mem[208][5] ),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(\cur_mb_mem[127][5] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(\cur_mb_mem[50][2] ),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(\cur_mb_mem[115][6] ),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(\best_cand_x[1] ),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(\cur_mb_mem[143][0] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(\min_sad_reg[6] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(\cur_mb_mem[68][1] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(\cur_mb_mem[153][4] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(\best_cand_x[3] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(\cur_mb_mem[24][0] ),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(\cur_mb_mem[224][4] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(\cur_mb_mem[140][0] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(\cur_mb_mem[192][4] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(\cur_mb_mem[91][1] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(\cur_mb_mem[45][3] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(\cur_mb_mem[134][6] ),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(\cur_mb_mem[150][6] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(\cur_mb_mem[50][0] ),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(\cur_mb_mem[85][0] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(\cur_mb_mem[164][1] ),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(\cur_mb_mem[28][2] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(\cur_mb_mem[151][3] ),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(\cur_mb_mem[41][1] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(\cur_mb_mem[88][6] ),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\cur_mb_mem[147][5] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(\cur_mb_mem[144][0] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(\cur_mb_mem[151][0] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(\cur_mb_mem[117][4] ),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(\cur_mb_mem[45][6] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(\cur_mb_mem[12][0] ),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(\cur_mb_mem[143][2] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(\cur_mb_mem[59][7] ),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(\cur_mb_mem[181][7] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(\cur_mb_mem[57][2] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(\cur_mb_mem[205][4] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(\cur_mb_mem[236][1] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(\cur_mb_mem[186][3] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(\cur_mb_mem[233][5] ),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(\cur_mb_mem[216][0] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(\cur_mb_mem[253][0] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(\cur_mb_mem[205][2] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(\cur_mb_mem[30][5] ),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(\cur_mb_mem[128][4] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(\cur_mb_mem[144][2] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(\current_accum_sad[8] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(\cur_mb_mem[252][7] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(\cur_mb_mem[47][7] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(\cur_mb_mem[157][2] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(\cur_mb_mem[144][3] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\cur_mb_mem[132][6] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(\cur_mb_mem[39][2] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\cur_mb_mem[157][4] ),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(\cur_mb_mem[188][2] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\cur_mb_mem[26][6] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(\cur_mb_mem[123][6] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\cur_mb_mem[177][7] ),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(\cur_mb_mem[185][0] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(\cur_mb_mem[182][1] ),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(\cur_mb_mem[136][6] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(\cur_mb_mem[221][2] ),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(\cur_mb_mem[249][6] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(\cur_mb_mem[1][4] ),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(\cur_mb_mem[245][7] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(\cur_mb_mem[29][0] ),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(\cur_mb_mem[236][7] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(\cur_mb_mem[230][0] ),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(\cur_mb_mem[213][3] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(\cur_mb_mem[245][6] ),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(\cur_mb_mem[4][5] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\cur_mb_mem[4][1] ),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(\cur_mb_mem[238][2] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(\cur_mb_mem[159][5] ),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(\cur_mb_mem[238][7] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(\cur_mb_mem[112][5] ),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(\cur_mb_mem[143][3] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(\cur_mb_mem[72][2] ),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(\cur_mb_mem[27][5] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(\cur_mb_mem[120][0] ),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(\cur_mb_mem[255][0] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(\cur_mb_mem[118][2] ),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(\cur_mb_mem[65][4] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(\cur_mb_mem[115][2] ),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(\cur_mb_mem[205][5] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(\cur_mb_mem[238][1] ),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(\cur_mb_mem[216][3] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(\cur_mb_mem[24][3] ),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(\cur_mb_mem[111][1] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(\cur_mb_mem[136][4] ),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(\cur_mb_mem[255][2] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(\cur_mb_mem[50][4] ),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(\cur_mb_mem[42][7] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\cur_mb_mem[134][2] ),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(\cur_mb_mem[128][3] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\cur_mb_mem[119][4] ),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(\cur_mb_mem[242][0] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(\cur_mb_mem[14][2] ),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(\cur_mb_mem[253][3] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(\cur_mb_mem[105][6] ),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(\cur_mb_mem[135][3] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(\cur_mb_mem[126][4] ),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(\cur_mb_mem[54][0] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(\cur_mb_mem[159][1] ),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(\cur_mb_mem[65][5] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(\cur_mb_mem[214][3] ),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(\cur_mb_mem[28][0] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(\cur_mb_mem[218][3] ),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(\cur_mb_mem[247][0] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(\cur_mb_mem[2][1] ),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(\cur_mb_mem[122][4] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(\cur_mb_mem[235][6] ),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(\cur_mb_mem[33][1] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(\cur_mb_mem[50][5] ),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(\cur_mb_mem[152][7] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(\cur_mb_mem[130][7] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(\cur_mb_mem[45][7] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(\cur_mb_mem[219][5] ),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(\cur_mb_mem[156][2] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(\cur_mb_mem[80][5] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(\cur_mb_mem[122][5] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\cur_mb_mem[193][1] ),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(\cur_mb_mem[226][4] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\cur_mb_mem[176][6] ),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(\cur_mb_mem[235][7] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(\cur_mb_mem[105][2] ),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(\cur_mb_mem[233][0] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(\cur_mb_mem[97][3] ),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(\cur_mb_mem[12][3] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(\cur_mb_mem[1][6] ),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(\cur_mb_mem[156][3] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(\cur_mb_mem[53][4] ),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(\cur_mb_mem[114][5] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(\cur_mb_mem[185][2] ),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(\cur_mb_mem[115][0] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(\cur_mb_mem[221][0] ),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(\cur_mb_mem[206][4] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(\cur_mb_mem[53][6] ),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(\cur_mb_mem[13][2] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(\cur_mb_mem[114][4] ),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(\cur_mb_mem[28][4] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(\cur_mb_mem[66][0] ),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(\cur_mb_mem[74][1] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(\cur_mb_mem[45][4] ),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(\cur_mb_mem[232][4] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(\cur_mb_mem[233][1] ),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(\cur_mb_mem[24][2] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(\cur_mb_mem[232][2] ),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(\cur_mb_mem[204][4] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(\cur_mb_mem[196][7] ),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(\cur_mb_mem[104][6] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(\cur_mb_mem[155][3] ),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(\cur_mb_mem[230][1] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(\cur_mb_mem[221][3] ),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(\cur_mb_mem[83][0] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(\cur_mb_mem[112][0] ),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(\cur_mb_mem[83][5] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(\cur_mb_mem[36][1] ),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(\cur_mb_mem[253][2] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(\cur_mb_mem[185][3] ),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(\cur_mb_mem[26][4] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(\cur_mb_mem[74][6] ),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(\cur_mb_mem[5][0] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(\cur_mb_mem[241][3] ),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(\cur_mb_mem[247][3] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(\cur_mb_mem[140][3] ),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(\cur_mb_mem[30][3] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(\cur_mb_mem[56][6] ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(\cur_mb_mem[30][2] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(\cur_mb_mem[242][5] ),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(\cur_mb_mem[246][3] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(\cur_mb_mem[226][5] ),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(\cur_mb_mem[200][3] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(\cur_mb_mem[232][3] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(\cur_mb_mem[80][4] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(\min_sad_reg[2] ),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(\cur_mb_mem[26][5] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(\cur_mb_mem[205][1] ),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(\cur_mb_mem[231][1] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(\cur_mb_mem[219][2] ),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(\cur_mb_mem[153][5] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(\cur_mb_mem[114][2] ),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(\min_sad_reg[5] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(\cur_mb_mem[177][0] ),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(\cur_mb_mem[67][4] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(\cur_mb_mem[11][6] ),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(\cur_mb_mem[153][1] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(\cur_mb_mem[119][5] ),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(\cur_mb_mem[5][2] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(\cur_mb_mem[154][1] ),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(\cur_mb_mem[52][6] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(\cur_mb_mem[37][2] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(\cur_mb_mem[180][7] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(\cur_mb_mem[238][6] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(\state[0] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(\best_cand_x[4] ),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(\cur_mb_mem[27][0] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\cur_mb_mem[97][0] ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(\cur_mb_mem[50][6] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\cur_mb_mem[45][5] ),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(\cur_mb_mem[129][6] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(\cur_mb_mem[120][1] ),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(\cur_mb_mem[5][3] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(\cur_mb_mem[241][4] ),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(\cur_mb_mem[240][5] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(\cur_mb_mem[200][5] ),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(\cur_mb_mem[234][3] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(\cur_mb_mem[31][3] ),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(\cur_mb_mem[97][6] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(\cur_mb_mem[112][2] ),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(\cur_mb_mem[10][3] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(\cur_mb_mem[29][2] ),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(\cur_mb_mem[204][5] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(\cur_mb_mem[233][3] ),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(\cur_mb_mem[65][6] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(\cur_mb_mem[148][2] ),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(\cur_mb_mem[209][1] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(\cur_mb_mem[242][4] ),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(\cur_mb_mem[209][5] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(\cur_mb_mem[35][2] ),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(\cur_mb_mem[240][4] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(\cur_mb_mem[206][5] ),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(\cur_mb_mem[142][6] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(\cur_mb_mem[135][7] ),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(\cur_mb_mem[142][7] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(\cur_mb_mem[247][2] ),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(\cur_mb_mem[0][6] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(net194),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(\cur_mb_mem[155][0] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(\cur_mb_mem[232][1] ),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(\cur_mb_mem[237][2] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\cur_mb_mem[231][4] ),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(\cur_mb_mem[236][6] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(\cur_mb_mem[120][2] ),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(\cur_mb_mem[148][3] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(\cur_mb_mem[206][1] ),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(\cur_mb_mem[25][1] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(net197),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(\cur_mb_mem[250][6] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(\cur_mb_mem[72][0] ),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(\min_sad_reg[9] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(\cur_mb_mem[83][1] ),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(\cur_mb_mem[31][5] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(\cur_mb_mem[108][0] ),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(\cur_mb_mem[233][2] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(\cur_mb_mem[228][2] ),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(\cur_mb_mem[11][1] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(\best_cand_x[2] ),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(\cur_mb_mem[240][1] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(\cur_mb_mem[232][5] ),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(\cur_mb_mem[23][6] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(\cur_mb_mem[124][3] ),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(\cur_mb_mem[241][5] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(\best_cand_x[5] ),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(\cur_mb_mem[234][5] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(\cur_mb_mem[120][3] ),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(\cur_mb_mem[135][2] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(\cur_mb_mem[108][3] ),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(\cur_mb_mem[209][7] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(\cur_mb_mem[151][2] ),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(\cur_mb_mem[102][6] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(\cur_mb_mem[120][5] ),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(\cur_mb_mem[12][2] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(\cur_mb_mem[148][0] ),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(\cur_mb_mem[228][5] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(\cur_mb_mem[236][2] ),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(\cur_mb_mem[138][6] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(\cur_mb_mem[214][2] ),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(\cur_mb_mem[131][7] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(\cur_mb_mem[177][3] ),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(\cur_mb_mem[135][0] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(\cur_mb_mem[108][2] ),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(\cur_mb_mem[128][1] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(\cur_mb_mem[84][2] ),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(\cur_mb_mem[219][0] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(\cur_mb_mem[146][7] ),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(\cur_mb_mem[207][2] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(\cur_mb_mem[219][3] ),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(\cur_mb_mem[83][4] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(\cur_mb_mem[234][6] ),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(\cur_mb_mem[195][5] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(\cur_mb_mem[26][2] ),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(\cur_mb_mem[213][7] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(\cur_mb_mem[235][5] ),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(\cur_mb_mem[236][3] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(\cur_mb_mem[195][4] ),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(\cur_mb_mem[158][7] ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(\cur_mb_mem[156][0] ),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(\best_cand_y[4] ),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(\cur_mb_mem[234][0] ),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(\cur_mb_mem[245][4] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(\cur_mb_mem[201][4] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(\cur_mb_mem[100][5] ),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(\cur_mb_mem[151][6] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(\cur_mb_mem[227][6] ),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(\cur_mb_mem[234][1] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(\cur_mb_mem[126][5] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(\cur_mb_mem[214][0] ),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(\cur_mb_mem[79][4] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(net193),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(\cur_mb_mem[88][0] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(\cur_mb_mem[238][0] ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(\cur_mb_mem[243][1] ),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(\cur_mb_mem[32][5] ),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(\cur_mb_mem[228][3] ),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(\cur_mb_mem[120][4] ),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(\cur_mb_mem[238][3] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(\cur_mb_mem[13][3] ),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(\cur_mb_mem[126][7] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(\cur_mb_mem[217][2] ),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(\cur_mb_mem[168][5] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(\cur_mb_mem[31][4] ),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(\cur_mb_mem[107][7] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(\cur_mb_mem[247][7] ),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(\cur_mb_mem[27][6] ),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(\cur_mb_mem[234][4] ),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(\cur_mb_mem[235][4] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(\cur_mb_mem[77][2] ),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(\cur_mb_mem[39][7] ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\cur_mb_mem[96][5] ),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(\cur_mb_mem[237][6] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(\cur_mb_mem[96][2] ),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(\cur_mb_mem[239][2] ),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(\cur_mb_mem[224][3] ),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(\shex_center_y[1] ),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(\cur_mb_mem[212][0] ),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(\cur_mb_mem[222][4] ),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(\cur_mb_mem[227][1] ),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(\cur_mb_mem[228][4] ),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(\shex_center_x[3] ),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(\cur_mb_mem[70][4] ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(\cur_mb_mem[201][5] ),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(\cur_mb_mem[222][5] ),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(\cur_mb_mem[33][6] ),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(\cur_mb_mem[29][3] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(\cur_mb_mem[230][3] ),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(\cur_mb_mem[32][4] ),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(\shex_center_x[6] ),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(\cur_mb_mem[13][0] ),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(\cur_mb_mem[237][3] ),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(\cur_mb_mem[129][7] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(\cur_mb_mem[69][4] ),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(\min_sad_reg[0] ),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(\cur_mb_mem[209][4] ),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(\cur_mb_mem[25][2] ),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(\shex_center_y[2] ),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(net184),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\cur_mb_mem[218][4] ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(\cur_mb_mem[255][3] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(\cur_mb_mem[221][5] ),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(\cur_mb_mem[155][7] ),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(\cur_mb_mem[131][3] ),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(\cur_mb_mem[104][2] ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\cur_mb_mem[198][0] ),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(\cur_mb_mem[30][6] ),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(\cur_mb_mem[128][7] ),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(\shex_center_y[3] ),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(\cur_mb_mem[97][2] ),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(\cur_mb_mem[104][0] ),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(\cur_mb_mem[214][4] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(\shex_center_x[5] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(\cur_mb_mem[96][0] ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(\cur_mb_mem[96][4] ),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(\cur_mb_mem[213][4] ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(\cur_mb_mem[213][5] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\cur_mb_mem[221][4] ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(\cur_mb_mem[202][2] ),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(\cur_mb_mem[70][7] ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(\shex_center_x[4] ),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(\shex_center_x[0] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(\min_sad_reg[15] ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(\cur_mb_mem[51][7] ),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(\cur_mb_mem[204][6] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(\cur_mb_mem[214][5] ),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(\cur_mb_mem[202][4] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(\cur_mb_mem[244][0] ),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(\cur_mb_mem[69][5] ),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(shex_load),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(\cur_mb_mem[218][5] ),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(\shex_center_y[6] ),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(\cur_mb_mem[54][6] ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(\min_sad_reg[1] ),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(\cur_mb_mem[248][3] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(\cur_mb_mem[123][4] ),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(\cur_mb_mem[54][2] ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\cur_mb_mem[203][4] ),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(\cur_mb_mem[5][1] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(\cur_mb_mem[100][4] ),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(\cur_mb_mem[4][3] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(\cur_mb_mem[198][5] ),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(\cur_mb_mem[232][0] ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(\cur_mb_mem[116][2] ),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(\cur_mb_mem[240][3] ),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(\cur_mb_mem[197][5] ),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(\cur_mb_mem[73][2] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(\cur_mb_mem[31][2] ),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(\cur_mb_mem[224][2] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\cur_mb_mem[245][3] ),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(\cur_mb_mem[215][7] ),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\cur_mb_mem[204][0] ),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(\cur_mb_mem[32][3] ),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\cur_mb_mem[197][4] ),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(\cur_mb_mem[38][7] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(\cur_mb_mem[131][0] ),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(\cand_x[3] ),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\state[0] ),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(\best_cand_y[1] ),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(\best_cand_y[1] ),
    .X(net1999));
 sky130_fd_sc_hd__buf_1 wire1 (.A(_08067_),
    .X(net2000));
 sky130_fd_sc_hd__clkbuf_1 max_cap2 (.A(net2002),
    .X(net2001));
 sky130_fd_sc_hd__clkbuf_1 wire3 (.A(_04819_),
    .X(net2002));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4 (.A(_06021_),
    .X(net2003));
 sky130_fd_sc_hd__clkbuf_1 max_cap5 (.A(_06004_),
    .X(net2004));
 sky130_fd_sc_hd__buf_1 wire6 (.A(_05992_),
    .X(net2005));
 sky130_fd_sc_hd__buf_1 max_cap7 (.A(_05974_),
    .X(net2006));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap8 (.A(_05894_),
    .X(net2007));
 sky130_fd_sc_hd__buf_1 wire9 (.A(_05889_),
    .X(net2008));
endmodule
